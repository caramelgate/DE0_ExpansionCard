DIGILENT
http://www.digilentinc.com/

PmodPS2 - Keyboard/mouse connector
http://www.digilentinc.com/Products/Detail.cfm?NavPath=2,401,529&Prod=PMOD-PS2
