

<!-- pf_header_start -->

<html>
  <head>
    <META NAME="keywords" CONTENT="cores, VHDL, Verilog HDL, ASIC, Synthesizable,
      standard cell, IP, Intellectual Property, 32-bit RISC, UART, PCI, SDRAM,
      full custom, system on a chip, SOC, reusable, design, development, synthesis,
      designs, developers, C, Linux, eCos, open, free, open source cores, RTL code,
      system-on-a-chip, circuits, digital, GNU, GPL, core, controller, processor,
      system design, chip design, EDA, design methodology, design tools, ASICs, programmable logic,
      FPGA's, PLDs, CPLDs, verification, Synthesis, HDL, Simulation, IC design software,
      semiconductor design, integrated circuits, system designs, chip designs, EDAs, 
      design methodologies, design tool, ASIC, programmable logics, FPGA, PLD, CPLD, Synthesis, 
      circuit, Synopsys, system design, chip design, programmable logic, FPGA's, PLDs, 
      CPLDs, verification, Simulation">
    <META NAME="description" CONTENT="OPENCORES.ORG endorses development and hosts
      a repository of free, open-source cores (chip designs) and supplemental
      platforms (boards).">
    <STYLE type=text/css>
      BODY {margin: 0;}
      BODY, P, DIV, TD, TR, TH, FORM, OL, UL, LI, B, I, INPUT, TEXTAREA, SELECT,
      FONT {font-size: 10pt; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}

      P, TD, FORM, TEXTAREA {font-size: 10pt;}

      H1, H2 {FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica; font-size: 13pt; text-decoration: none}

      .noline {text-decoration: none;}

      .menu_top {text-decoration: none; font-weight: bold;
        font-size: 7pt; color: #000000; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;} 
      .menu_section {text-decoration: none; font-weight: bold;
        font-size: 10pt; color: #ffffff; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;} 
      .menu_item {font-size: 10pt; color: #004488; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}
      .menu_section_admin {text-decoration: none; font-weight: bold;
        font-size: 10pt; color: #ffff44; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;} 
      .page_title {text-decoration: none; font-weight: bold; color: #c00000; font-size: 13pt; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}
      .block_title {text-decoration: none; font-weight: bold; font-size: 11pt; color: #000000; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}
      .block_subtitle {text-decoration: none; font-weight: bold; font-size: 10pt; color: #000000; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}
      .title {text-decoration: none; font-weight: bold; font-size: 10pt; color: #000000; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}

      .large {font-size: 13pt; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}
      .medium {font-size: 10pt; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}
      .small {font-size: 7pt; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}
      .ultrasmall {font-size: 3pt; FONT-FAMILY: Verdana, Tahoma, Arial, Helvetica;}

      .button { font-family:Verdana, Tahoma, Arial, Helvetica; }
      .searchfield {font-family: verdana, arial, helvetica; font-size: 10px; color: #333333; width: 80px; height: 17px;}

    </STYLE>

    <title>OPENCORES.ORG</title>

    <script laguage="Javascript">
      function check(msg) {
        if(confirm(msg)) {
          return true
        } else {
          return false
        }
      }
    </script>

<script src="http://www.google-analytics.com/urchin.js"
type="text/javascript">

</script>

<script type="text/javascript">

_uacct = "UA-2763846-2";

urchinTracker();

</script>

  </head>

  

  <body 
    bgcolor="#e0e0e0" 
    topmargin="0" 
    leftmargin="0" 
    marginwidth="0" 
    marginheight="0" 
    link="#004488" 
    alink="#ff3300"
    vlink="#444444"
  >

<a name="top">
<!-- pf_header_end -->
<center>
<table cellpadding=0 cellspacing=0 border=0 width=96%><tr>
<td width=1 bgcolor=#000000><img width=1 src="/images/dotty.gif"></td>

<td>

<table border=0 cellpadding=0 cellspacing=0 width=100%>

<tr><td bgcolor="#ffffff" height=70>

<table width=100% border=0 ><tr>
<td valign=center width="30"><img height=1 width=30 src="/images/dotty.gif"></td>
<td width=70 valign=center>
<a href="/"><img style="padding-left: 0px;" border=0 src="/images/newlogo.gif"></a>
</td><td>
<a href="/"><img style="padding-left: 0px;"  align=baseline border=0 src="/images/newlogotext.gif"></a>
</td><td>
<center>

<!--
<a title="" href="/banner.cgi/redirect/14"><img width=468 height=60 border=0 alt="" src="/banner.cgi/iframe/14"></a>
//-->

</center>
</td><td align=right>


<iframe frameborder=0 scrolling=0 marginwidth=0 marignheight=0 width=304 height=63
  leftmargin="0" topmargin="0" hspace=0 vspace=0 src="http://www.opencores.org/banner.cgi/iframe/14"></iframe>






</td>
</tr></table>

</td></tr>
<tr bgcolor=#000000><td><img height=1 src="/images/dotty.gif"></td></tr>
<tr><td bgcolor=#ffffff>


<table border=0 cellpadding=0 cellspacing=0 width=100%><tr>

<td bgcolor=#b3b3b3 width=60% background="/images/menu1.gif"></td>
<td bgcolor=#b3b3b3 width=15 background="/images/menu1.gif" align=right><img border=0 src="/images/exp1.gif"></td>

<td bgcolor=#ffffff align=right nowrap>
&nbsp; &nbsp; &nbsp; &nbsp; 
<font class=menu_top size=-1>
        
          <a class=menu_top href="/login.cgi/login">LOGIN</a>
          
            &nbsp; ::: &nbsp;
          
        
          <a class=menu_top href="/recover_pass.cgi/recover_pass">RECOVER PASS</a>
          
            &nbsp; ::: &nbsp;
          
        
          <a class=menu_top href="/get_account.cgi/get_account">FOR DEVELOPERS</a>
          
        

&nbsp; &nbsp;
</font>

</td></tr>
<tr bgcolor=#ffffff>
  <td></td>
  <td></td>
  <td bgcolor=#000000><img src="/images/dotty.gif"></td>
</tr>

</table>

<table border=0 cellpadding=0 cellspacing=0>
<tr>
<td width=10><img width=10 src="/images/dotty.gif"></td>

<td width=120 valign=top>
        
        <table width=100% border=0 cellpadding=2 cellspacing=0>
          <tr><td><img height=2 src="/images/dotty.gif"></td></tr>
        
         <tr><td bgcolor="#347FB8">
           <img src="/images/bullet.gif">
         
           <font class=menu_section>Browse</font>
         
         </td></tr>
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/browse.cgi/by_category"><font class=menu_item>Projects</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/cvsweb.shtml/"><font class=menu_item>Code (CVS)</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/forums.cgi"><font class=menu_item>Forums</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/news.cgi/list/1"><font class=menu_item>News</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/articles.cgi/list"><font class=menu_item>Articles</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/polls.cgi/list"><font class=menu_item>Polls</font></a></li>
            
           </td></tr>
            
          
          <tr><td><font size=-2>&nbsp;</font></td></tr>
        
         <tr><td bgcolor="#347FB8">
           <img src="/images/bullet.gif">
         
           <font class=menu_section>OpenCores</font>
         
         </td></tr>
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/faq.cgi/index"><font class=menu_item>FAQ</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/cvs_howto"><font class=menu_item>CVS HowTo</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/mission"><font class=menu_item>Mission</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/media"><font class=menu_item>Media</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/tools"><font class=menu_item>Tools</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/sponsors"><font class=menu_item>Sponsors</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/mirrors"><font class=menu_item>Mirrors</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/logos"><font class=menu_item>Logos</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opencores/contacts"><font class=menu_item>Contact us</font></a></li>
            
           </td></tr>
            
          
          <tr><td><font size=-2>&nbsp;</font></td></tr>
        
         <tr><td bgcolor="#347FB8">
           <img src="/images/bullet.gif">
         
           <font class=menu_section>Tools</font>
         
         </td></tr>
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <font class=menu_item><a href="/search.cgi">Search</a><br><table><tr><form action=/search.cgi/do_search><td><font class=small>&nbsp;&nbsp;</font></td><td><input class=searchfield type=text name=query></td></form></tr></table></font></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/cvsget.shtml"><font class=menu_item>Download Cores (CVSGet)</font></a></li>
            
           </td></tr>
            
          
          <tr><td><font size=-2>&nbsp;</font></td></tr>
        
         <tr><td bgcolor="#347FB8">
           <img src="/images/bullet.gif">
         
           <font class=menu_section>More</font>
         
         </td></tr>
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/wishbone/"><font class=menu_item>Wishbone</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/perlilog/"><font class=menu_item>Perlilog</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/edatools/"><font class=menu_item>EDA tools</font></a></li>
            
           </td></tr>
            
          
           <tr><td>
              
                  
                      <li class=small>
                  
              
            
                <a class=menu_item href="/projects.cgi/web/opentech/"><font class=menu_item>OpenTech CD</font></a></li>
            
           </td></tr>
            
          
          <tr><td><font size=-2>&nbsp;</font></td></tr>
        
        </table>



</td>
<td width=10><img width=10 src="/images/dotty.gif"></td>
<td background="/images/vpd.gif"><img width=1 src="/images/dotty.gif"></td>
<td width=10><img width=10 src="/images/dotty.gif"></td>
<td valign=top>


        
        <table width=100% cellpadding=2 cellspacing=0 border=0>
          <tr><td><img height=2 src="/images/dotty.gif"></td></tr>
        </table>
        


<table width=100% cellspacing=0 cellpadding=0 border=0><tr><td>

<!-- pf_body_start -->







 

<!DOCTYPE html PUBLIC "-//W3C//DTD XHTML 1.0 Transitional//EN" "http://www.w3.org/TR/xhtml1/DTD/xhtml1-transitional.dtd">
<html>
<head>
<title>CVS log for spdif_interface/rtl/vhdl/tx_bitbuf.vhd</title>
<meta name="robots" content="nofollow" />
<meta name="generator" content="FreeBSD-CVSweb 3.0.5" />
<meta http-equiv="Content-Script-Type" content="text/javascript" />
<meta http-equiv="Content-Style-Type" content="text/css" />
<link rel="stylesheet" type="text/css" href="/css/cvsweb.css" />
</head>
<body>
 <h1>CVS log for spdif_interface/rtl/vhdl/tx_bitbuf.vhd</h1>
<p>
 <a href="./#tx_bitbuf.vhd"><img src="/icons/back.gif" alt="[BACK]" border="0" width="20" height="22" /></a> <b>Up to  <a href="/cvsweb.shtml/#dirlist">[Official OpenCores CVS Repository]</a> / <a href="/cvsweb.shtml/spdif_interface/#dirlist">spdif_interface</a> / <a href="/cvsweb.shtml/spdif_interface/rtl/#dirlist">rtl</a> / <a href="/cvsweb.shtml/spdif_interface/rtl/vhdl/#dirlist">vhdl</a></b>
</p>
<p>
 <a href="#diff">Request diff between arbitrary revisions</a>
</p>
<hr />
<p>
Keyword substitution: kv<br />
Default branch: MAIN<br />
</p>
<hr />
<a name="rev1.4"></a><a name="HEAD"></a><a name="MAIN"></a>
 Revision <b>1.4</b>: <a href="/cvsweb.cgi/~checkout~/spdif_interface/rtl/vhdl/tx_bitbuf.vhd?rev=1.4;content-type=text%2Fplain" class="download-link">download</a> - view: <a href="tx_bitbuf.vhd?rev=1.4;content-type=text%2Fplain" class="display-link">text</a>, <a href="tx_bitbuf.vhd?rev=1.4;content-type=text%2Fx-cvsweb-markup" class="display-link">markup</a>, <a href="tx_bitbuf.vhd?annotate=1.4">annotated</a> - <a href="tx_bitbuf.vhd?r1=1.4#rev1.4">select&nbsp;for&nbsp;diffs</a><br />
<i>Thu Oct 11 19:14:43 2007 UTC</i> (3 months, 2 weeks ago) by <i>gedra</i><br />
Branches: <a href="./tx_bitbuf.vhd?only_with_tag=MAIN">MAIN</a><br />
CVS tags: <a href="./tx_bitbuf.vhd?only_with_tag=HEAD">HEAD</a><br />
Diff to previous 1.3: <a href="tx_bitbuf.vhd.diff?r1=1.3;r2=1.4">preferred</a>, <a href="tx_bitbuf.vhd.diff?r1=1.3;r2=1.4;f=u">unified</a><br />
Changes since revision 1.3: +45 -42 lines<br />
<pre class="log">
Code beautification
</pre>
<hr />
<a name="rev1.3"></a><a name="spdif_rel_1"></a><a name="beta_2"></a>
 Revision <b>1.3</b>: <a href="/cvsweb.cgi/~checkout~/spdif_interface/rtl/vhdl/tx_bitbuf.vhd?rev=1.3;content-type=text%2Fplain" class="download-link">download</a> - view: <a href="tx_bitbuf.vhd?rev=1.3;content-type=text%2Fplain" class="display-link">text</a>, <a href="tx_bitbuf.vhd?rev=1.3;content-type=text%2Fx-cvsweb-markup" class="display-link">markup</a>, <a href="tx_bitbuf.vhd?annotate=1.3">annotated</a> - <a href="tx_bitbuf.vhd?r1=1.3#rev1.3">select&nbsp;for&nbsp;diffs</a><br />
<i>Mon Jul 19 16:59:43 2004 UTC</i> (3 years, 6 months ago) by <i>gedra</i><br />
Branches: <a href="./tx_bitbuf.vhd?only_with_tag=MAIN">MAIN</a><br />
CVS tags: <a href="./tx_bitbuf.vhd?only_with_tag=spdif_rel_1">spdif_rel_1</a>,
<a href="./tx_bitbuf.vhd?only_with_tag=beta_2">beta_2</a><br />
Diff to previous 1.2: <a href="tx_bitbuf.vhd.diff?r1=1.2;r2=1.3">preferred</a>, <a href="tx_bitbuf.vhd.diff?r1=1.2;r2=1.3;f=u">unified</a><br />
Changes since revision 1.2: +16 -6
 lines<br />
<pre class="log">
Fixed bug.
</pre>
<hr />
<a name="rev1.2"></a>
 Revision <b>1.2</b>: <a href="/cvsweb.cgi/~checkout~/spdif_interface/rtl/vhdl/tx_bitbuf.vhd?rev=1.2;content-type=text%2Fplain" class="download-link">download</a> - view: <a href="tx_bitbuf.vhd?rev=1.2;content-type=text%2Fplain" class="display-link">text</a>, <a href="tx_bitbuf.vhd?rev=1.2;content-type=text%2Fx-cvsweb-markup" class="display-link">markup</a>, <a href="tx_bitbuf.vhd?annotate=1.2">annotated</a> - <a href="tx_bitbuf.vhd?r1=1.2#rev1.2">select&nbsp;for&nbsp;diffs</a><br />
<i>Sat Jul 17 17:21:11 2004 UTC</i> (3 years, 6 months ago) by <i>gedra</i><br />
Branches: <a href="./tx_bitbuf.vhd?only_with_tag=MAIN">MAIN</a><br />
Diff to previous 1.1: <a href="tx_bitbuf.vhd.diff?r1=1.1;r2=1.2">preferred</a>, <a href="tx_bitbuf.vhd.diff?r1=1.1;r2=1.2;f=u">unified</a><br />
Changes since revision 1.1: +6 -3
 lines<br />
<pre class="log">
Fixed bug.
</pre>
<hr />
<a name="rev1.1"></a>
 Revision <b>1.1</b>: <a href="/cvsweb.cgi/~checkout~/spdif_interface/rtl/vhdl/tx_bitbuf.vhd?rev=1.1;content-type=text%2Fplain" class="download-link">download</a> - view: <a href="tx_bitbuf.vhd?rev=1.1;content-type=text%2Fplain" class="display-link">text</a>, <a href="tx_bitbuf.vhd?rev=1.1;content-type=text%2Fx-cvsweb-markup" class="display-link">markup</a>, <a href="tx_bitbuf.vhd?annotate=1.1">annotated</a> - <a href="tx_bitbuf.vhd?r1=1.1#rev1.1">select&nbsp;for&nbsp;diffs</a><br />
<i>Wed Jul 14 17:58:19 2004 UTC</i> (3 years, 6 months ago) by <i>gedra</i><br />
Branches: <a href="./tx_bitbuf.vhd?only_with_tag=MAIN">MAIN</a><br />
<pre class="log">
Transmitter channel status buffer.
</pre>
<hr />
<form method="get" action="/cvsweb.shtml/spdif_interface/rtl/vhdl/tx_bitbuf.vhd.diff" id="diff_select">
<fieldset>
<legend>Diff request</legend>
<p>
 <a name="diff">
  This form allows you to request diffs between any two revisions of a file.
  You may select a symbolic revision name using the selection box or you may
  type in a numeric name using the type-in text box.
 </a>
</p>
<table summary="Diff between arbitrary revisions">
<tr>
<td class="opt-label">
<label for="r1" accesskey="1">Diffs between</label>
</td>
<td class="opt-value">
<select id="r1" name="r1">
<option value="text" selected="selected">Use Text Field</option>
<option value="1.3:spdif_rel_1">spdif_rel_1</option>
<option value="1.3:beta_2">beta_2</option>
<option value="1:MAIN">MAIN</option>
<option value="1.4:HEAD">HEAD</option>
</select>
<input type="text" size="12" name="tr1" value="1.1" onchange="this.form.r1.selectedIndex=0" />
</td>
<td></td>
</tr>
<tr>
<td class="opt-label">
<label for="r2" accesskey="2">and</label>
</td>
<td class="opt-value">
<select id="r2" name="r2">
<option value="text" selected="selected">Use Text Field</option>
<option value="1.3:spdif_rel_1">spdif_rel_1</option>
<option value="1.3:beta_2">beta_2</option>
<option value="1:MAIN">MAIN</option>
<option value="1.4:HEAD">HEAD</option>
</select>
<input type="text" size="12" name="tr2" value="1.4" onchange="this.form.r2.selectedIndex=0" />
</td>
<td><input type="submit" value="Get Diffs" accesskey="G" /></td>
</tr>
</table>
</fieldset>
</form>
<form method="get" action="/cvsweb.shtml/spdif_interface/rtl/vhdl/tx_bitbuf.vhd">
<fieldset>
<legend>Log view options</legend>
<table summary="Log view options">
<tr>
<td class="opt-label">
<label for="f" accesskey="D">Preferred diff type:</label>
</td>
<td class="opt-value">
<select id="f" name="f" onchange="this.form.submit()">
<option value="h" selected="selected">Colored</option>
<option value="H">Long colored</option>
<option value="u">Unified</option>
<option value="c">Context</option>
<option value="s">Side by side</option>
</select></td>
<td></td>
</tr>
<tr>
<td class="opt-label">
<label for="only_with_tag" accesskey="B">View only branch:</label>
</td>
<td class="opt-value">
<a name="branch">
<select id="only_with_tag" name="only_with_tag" onchange="this.form.submit()">
<option value="" selected="selected">Show all branches</option>
<option>MAIN</option></select>
</a>
</td>
<td></td>
</tr>
<tr>
<td class="opt-label">
<label for="logsort" accesskey="L">Sort log by:</label>
</td>
<td>
<select id="logsort" name="logsort" onchange="this.form.submit()">
<option value="cvs">Not sorted</option>
<option value="date" selected="selected">Commit date</option>
<option value="rev">Revision</option>
</select></td>
<td><input type="submit" value="Set" accesskey="S" /></td>
</tr>
</table>
</fieldset>
</form>
<hr />
<address><span style="font-size: smaller">FreeBSD-CVSweb &lt;<a href="mailto:freebsd-cvsweb@FreeBSD.org">freebsd-cvsweb@FreeBSD.org</a>&gt;</span></address>
</body>
</html>







<!-- pf_body_end -->

</td>
<td><img width=15 src="/images/dotty.gif"></td>
</tr></table>

<xcenter>

<img border=0 src="/images/dotty.gif" height=1 width=400>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>
<img border=0 src="/images/dotty.gif" height=1 width=30>

</td></tr>
</table>

&nbsp;

</td></tr>

<tr bgcolor=#000000><td><img height=1 src="/images/dotty.gif"></td></tr>
</table>

<table bgcolor="b3b3b3" width=100% cellpadding=0 cellspacing=0 border=0>
<tr><td align=right>
Copyright (c) 1999-2007 OPENCORES.ORG. All rights reserved. &nbsp;
</td></tr>
<tr><td>
&nbsp;
</td></tr>
</table>

</td>
<td width=1 bgcolor=#000000><img width=1 src="/images/dotty.gif"></td>
<td width=1 bgcolor=#f0f0c8><img width=1 src="/images/dotty.gif"></td>
</tr></table>
</center>

<!-- pf_footer_start -->

  </body>
</html>

<!-- pf_footer_end -->



