// megafunction wizard: %ALTLVDS%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altlvds_tx 

// ============================================================
// File Name: alt_diff_out_x4_raw.v
// Megafunction Name(s):
// 			altlvds_tx
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module alt_diff_out_x4_raw (
	tx_in,
	tx_inclock,
	tx_syncclock,
	tx_out);

	input	[39:0]  tx_in;
	input	  tx_inclock;
	input	  tx_syncclock;
	output	[3:0]  tx_out;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	  tx_syncclock;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [3:0] sub_wire0;
	wire [3:0] tx_out = sub_wire0[3:0];

	altlvds_tx	altlvds_tx_component (
				.tx_in (tx_in),
				.tx_syncclock (tx_syncclock),
				.tx_inclock (tx_inclock),
				.tx_out (sub_wire0),
				.pll_areset (1'b0),
				.sync_inclock (1'b0),
				.tx_coreclock (),
				.tx_data_reset (1'b0),
				.tx_enable (1'b1),
				.tx_locked (),
				.tx_outclock (),
				.tx_pll_enable (1'b1));
	defparam
		altlvds_tx_component.deserialization_factor = 10,
		altlvds_tx_component.implement_in_les = "ON",
		altlvds_tx_component.intended_device_family = "Cyclone III",
		altlvds_tx_component.lpm_hint = "CBX_MODULE_PREFIX=alt_diff_out_x4_raw",
		altlvds_tx_component.lpm_type = "altlvds_tx",
		altlvds_tx_component.number_of_channels = 4,
		altlvds_tx_component.registered_input = "OFF",
		altlvds_tx_component.use_external_pll = "ON";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: Deser_Factor NUMERIC "10"
// Retrieval info: PRIVATE: Enable_DPA_Mode STRING "OFF"
// Retrieval info: PRIVATE: Ext_PLL STRING "ON"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: Int_Device STRING "Cyclone III"
// Retrieval info: PRIVATE: LVDS_Mode NUMERIC "0"
// Retrieval info: PRIVATE: Le_Serdes STRING "ON"
// Retrieval info: PRIVATE: Num_Channel NUMERIC "4"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "10"
// Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "ON"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_tx"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "4"
// Retrieval info: CONSTANT: REGISTERED_INPUT STRING "OFF"
// Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "ON"
// Retrieval info: USED_PORT: tx_in 0 0 40 0 INPUT NODEFVAL tx_in[39..0]
// Retrieval info: USED_PORT: tx_inclock 0 0 0 0 INPUT_CLK_EXT GND tx_inclock
// Retrieval info: USED_PORT: tx_out 0 0 4 0 OUTPUT NODEFVAL tx_out[3..0]
// Retrieval info: USED_PORT: tx_syncclock 0 0 0 0 INPUT GND tx_syncclock
// Retrieval info: CONNECT: @tx_in 0 0 40 0 tx_in 0 0 40 0
// Retrieval info: CONNECT: tx_out 0 0 4 0 @tx_out 0 0 4 0
// Retrieval info: CONNECT: @tx_syncclock 0 0 0 0 tx_syncclock 0 0 0 0
// Retrieval info: CONNECT: @tx_inclock 0 0 0 0 tx_inclock 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_diff_out_x4_raw.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_diff_out_x4_raw.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_diff_out_x4_raw.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_diff_out_x4_raw.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_diff_out_x4_raw.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_diff_out_x4_raw_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_diff_out_x4_raw_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
// Retrieval info: CBX_MODULE_PREFIX: ON
