//
// 16Bit x 4K synched ROM
//
module sub_rom(
  CLK,
  A,
  DO
);

input  CLK;
input  [10:0] A;
output [15:0] DO;

reg [15:0] DO;

function [15:0] rom ;
input [10:0] addr;
begin
case(addr)
  11'h0:rom=16'h112;
  11'h1:rom=16'h14;
  11'h2:rom=16'hA0;
  11'h3:rom=16'h624;
  11'h4:rom=16'hB16;
  11'h5:rom=16'hF21;
  11'h6:rom=16'hF11;
  11'h7:rom=16'hF01;
  11'h8:rom=16'hFF1;
  11'h9:rom=16'hF90;
  11'hA:rom=16'h1FF1;
  11'hB:rom=16'h8801;
  11'hC:rom=16'hC801;
  11'hD:rom=16'h2705;
  11'hE:rom=16'h29F2;
  11'hF:rom=16'hC802;
  11'h10:rom=16'h2107;
  11'h11:rom=16'hC804;
  11'h12:rom=16'h2110;
  11'h13:rom=16'hC808;
  11'h14:rom=16'h212A;
  11'h15:rom=16'hFF1;
  11'h16:rom=16'hF90;
  11'h17:rom=16'h1F01;
  11'h18:rom=16'hC07;
  11'h19:rom=16'h308D;
  11'h1A:rom=16'h29ED;
  11'h1B:rom=16'h27F4;
  11'h1C:rom=16'h8024;
  11'h1D:rom=16'h1C07;
  11'h1E:rom=16'hE01;
  11'h1F:rom=16'h6010;
  11'h20:rom=16'h1E01;
  11'h21:rom=16'h2FE6;
  11'h22:rom=16'h1F01;
  11'h23:rom=16'hC06;
  11'h24:rom=16'h9001;
  11'h25:rom=16'h23E2;
  11'h26:rom=16'h1C06;
  11'h27:rom=16'h29E0;
  11'h28:rom=16'hC05;
  11'h29:rom=16'hC080;
  11'h2A:rom=16'h2907;
  11'h2B:rom=16'hC040;
  11'h2C:rom=16'h290C;
  11'h2D:rom=16'h1F11;
  11'h2E:rom=16'h2704;
  11'h2F:rom=16'h2F53;
  11'h30:rom=16'h2FD6;
  11'h31:rom=16'h7002;
  11'h32:rom=16'h1E02;
  11'h33:rom=16'h70EA;
  11'h34:rom=16'h1C06;
  11'h35:rom=16'h7040;
  11'h36:rom=16'h1C05;
  11'h37:rom=16'h2FD0;
  11'h38:rom=16'h7003;
  11'h39:rom=16'h1E02;
  11'h3A:rom=16'h1F11;
  11'h3B:rom=16'h2704;
  11'h3C:rom=16'h2F53;
  11'h3D:rom=16'h2FC9;
  11'h3E:rom=16'h1F01;
  11'h3F:rom=16'h1F11;
  11'h40:rom=16'h1F21;
  11'h41:rom=16'h2711;
  11'h42:rom=16'h7200;
  11'h43:rom=16'h200;
  11'h44:rom=16'h211;
  11'h45:rom=16'h301D;
  11'h46:rom=16'h28BF;
  11'h47:rom=16'h10;
  11'h48:rom=16'hC201;
  11'h49:rom=16'h2103;
  11'h4A:rom=16'h2701;
  11'h4B:rom=16'hF100;
  11'h4C:rom=16'h1E1B;
  11'h4D:rom=16'h8001;
  11'h4E:rom=16'h1200;
  11'h4F:rom=16'h2FB6;
  11'h50:rom=16'h1FF1;
  11'h51:rom=16'h1F01;
  11'h52:rom=16'h1F11;
  11'h53:rom=16'hC05;
  11'h54:rom=16'hC0C0;
  11'h55:rom=16'h2923;
  11'h56:rom=16'hC04;
  11'h57:rom=16'h2780;
  11'h58:rom=16'hF000;
  11'h59:rom=16'hE12;
  11'h5A:rom=16'h4101;
  11'h5B:rom=16'h2103;
  11'h5C:rom=16'h2780;
  11'h5D:rom=16'h5000;
  11'h5E:rom=16'h1C04;
  11'h5F:rom=16'hC05;
  11'h60:rom=16'h9001;
  11'h61:rom=16'h1C05;
  11'h62:rom=16'h2104;
  11'h63:rom=16'h700F;
  11'h64:rom=16'h1C06;
  11'h65:rom=16'h2F0F;
  11'h66:rom=16'h1F21;
  11'h67:rom=16'h1F31;
  11'h68:rom=16'h1F41;
  11'h69:rom=16'h1F51;
  11'h6A:rom=16'h1F61;
  11'h6B:rom=16'h1F71;
  11'h6C:rom=16'h2702;
  11'h6D:rom=16'h2FD7;
  11'h6E:rom=16'hF71;
  11'h6F:rom=16'hF61;
  11'h70:rom=16'hF51;
  11'h71:rom=16'hF41;
  11'h72:rom=16'hF31;
  11'h73:rom=16'hF21;
  11'h74:rom=16'hF11;
  11'h75:rom=16'hF01;
  11'h76:rom=16'hFF1;
  11'h77:rom=16'hF90;
  11'h78:rom=16'hC080;
  11'h79:rom=16'h29FB;
  11'h7A:rom=16'hC04;
  11'h7B:rom=16'h7102;
  11'h7C:rom=16'hC001;
  11'h7D:rom=16'h2102;
  11'h7E:rom=16'h5101;
  11'h7F:rom=16'h1E12;
  11'h80:rom=16'hE12;
  11'h81:rom=16'h2780;
  11'h82:rom=16'hF000;
  11'h83:rom=16'h2904;
  11'h84:rom=16'h3017;
  11'h85:rom=16'h2704;
  11'h86:rom=16'h2F53;
  11'h87:rom=16'h1C04;
  11'h88:rom=16'h2FEC;
  11'h89:rom=16'h2718;
  11'h8A:rom=16'h7F00;
  11'h8B:rom=16'h2720;
  11'h8C:rom=16'h7E00;
  11'h8D:rom=16'h2710;
  11'h8E:rom=16'h7D80;
  11'h8F:rom=16'h2710;
  11'h90:rom=16'h7C92;
  11'h91:rom=16'h2710;
  11'h92:rom=16'h7B00;
  11'h93:rom=16'h2710;
  11'h94:rom=16'h7AD8;
  11'h95:rom=16'h7800;
  11'h96:rom=16'hE05;
  11'h97:rom=16'h7003;
  11'h98:rom=16'h1E02;
  11'h99:rom=16'h7000;
  11'h9A:rom=16'h1E01;
  11'h9B:rom=16'h7000;
  11'h9C:rom=16'h1E0D;
  11'h9D:rom=16'h2710;
  11'h9E:rom=16'h7000;
  11'h9F:rom=16'h2718;
  11'hA0:rom=16'h7100;
  11'hA1:rom=16'h7200;
  11'hA2:rom=16'h1020;
  11'hA3:rom=16'h8002;
  11'hA4:rom=16'h301D;
  11'hA5:rom=16'h29FD;
  11'hA6:rom=16'h270E;
  11'hA7:rom=16'h2F1F;
  11'hA8:rom=16'h2701;
  11'hA9:rom=16'h705E;
  11'hAA:rom=16'h7150;
  11'hAB:rom=16'h2718;
  11'hAC:rom=16'h7200;
  11'hAD:rom=16'h2705;
  11'hAE:rom=16'h2F7E;
  11'hAF:rom=16'h27FF;
  11'hB0:rom=16'h70F7;
  11'hB1:rom=16'h1C01;
  11'hB2:rom=16'h2710;
  11'hB3:rom=16'h70B8;
  11'hB4:rom=16'h71FF;
  11'hB5:rom=16'h1D01;
  11'hB6:rom=16'h1D02;
  11'hB7:rom=16'h1010;
  11'hB8:rom=16'h7001;
  11'hB9:rom=16'h71FF;
  11'hBA:rom=16'h1D04;
  11'hBB:rom=16'h1D15;
  11'hBC:rom=16'h7003;
  11'hBD:rom=16'h1C00;
  11'hBE:rom=16'h2702;
  11'hBF:rom=16'h2FCD;
  11'hC0:rom=16'h2706;
  11'hC1:rom=16'h703A;
  11'hC2:rom=16'h7150;
  11'hC3:rom=16'h7200;
  11'hC4:rom=16'h2705;
  11'hC5:rom=16'h2F8B;
  11'hC6:rom=16'h2701;
  11'hC7:rom=16'h7000;
  11'hC8:rom=16'h710E;
  11'hC9:rom=16'h1E0C;
  11'hCA:rom=16'h1E1D;
  11'hCB:rom=16'h70FF;
  11'hCC:rom=16'h2704;
  11'hCD:rom=16'h2F5D;
  11'hCE:rom=16'h3F90;
  11'hCF:rom=16'hE01;
  11'hD0:rom=16'hC002;
  11'hD1:rom=16'h2104;
  11'hD2:rom=16'h2701;
  11'hD3:rom=16'h2FB1;
  11'hD4:rom=16'h2FFB;
  11'hD5:rom=16'h2702;
  11'hD6:rom=16'h2F7F;
  11'hD7:rom=16'h2FF8;
  11'hD8:rom=16'h2710;
  11'hD9:rom=16'h7080;
  11'hDA:rom=16'h7101;
  11'hDB:rom=16'h2704;
  11'hDC:rom=16'h2FA9;
  11'hDD:rom=16'hD00;
  11'hDE:rom=16'hD0F0;
  11'hDF:rom=16'h2808;
  11'hE0:rom=16'hD0E0;
  11'hE1:rom=16'h281C;
  11'hE2:rom=16'hD0D8;
  11'hE3:rom=16'h2815;
  11'hE4:rom=16'hD0D0;
  11'hE5:rom=16'h280E;
  11'hE6:rom=16'hF00;
  11'hE7:rom=16'hD0F0;
  11'hE8:rom=16'h2102;
  11'hE9:rom=16'hF00;
  11'hEA:rom=16'h2710;
  11'hEB:rom=16'h70B6;
  11'hEC:rom=16'h7102;
  11'hED:rom=16'h2704;
  11'hEE:rom=16'h2FA9;
  11'hEF:rom=16'h9002;
  11'hF0:rom=16'h00;
  11'hF1:rom=16'h1E07;
  11'hF2:rom=16'hF00;
  11'hF3:rom=16'h2710;
  11'hF4:rom=16'h70A4;
  11'hF5:rom=16'h7106;
  11'hF6:rom=16'h2704;
  11'hF7:rom=16'h2FA8;
  11'hF8:rom=16'h2710;
  11'hF9:rom=16'h70A4;
  11'hFA:rom=16'h7106;
  11'hFB:rom=16'h2704;
  11'hFC:rom=16'h2FCA;
  11'hFD:rom=16'h400F;
  11'hFE:rom=16'hE004;
  11'hFF:rom=16'h2702;
  11'h100:rom=16'h800A;
  11'h101:rom=16'h20;
  11'h102:rom=16'h01;
  11'h103:rom=16'h7101;
  11'h104:rom=16'h3F22;
  11'h105:rom=16'h19E;
  11'h106:rom=16'h00;
  11'h107:rom=16'h19E;
  11'h108:rom=16'h00;
  11'h109:rom=16'h19E;
  11'h10A:rom=16'h00;
  11'h10B:rom=16'h24A;
  11'h10C:rom=16'h10B2;
  11'h10D:rom=16'h250;
  11'h10E:rom=16'h1086;
  11'h10F:rom=16'h19E;
  11'h110:rom=16'h00;
  11'h111:rom=16'h25A;
  11'h112:rom=16'h00;
  11'h113:rom=16'h262;
  11'h114:rom=16'h10A2;
  11'h115:rom=16'h4CA;
  11'h116:rom=16'h10A2;
  11'h117:rom=16'h268;
  11'h118:rom=16'h1088;
  11'h119:rom=16'h4CA;
  11'h11A:rom=16'h1088;
  11'h11B:rom=16'h4CA;
  11'h11C:rom=16'h108A;
  11'h11D:rom=16'h26E;
  11'h11E:rom=16'h10AA;
  11'h11F:rom=16'h24A;
  11'h120:rom=16'h10AA;
  11'h121:rom=16'h276;
  11'h122:rom=16'h10AE;
  11'h123:rom=16'h24A;
  11'h124:rom=16'h10AE;
  11'h125:rom=16'h7103;
  11'h126:rom=16'h2704;
  11'h127:rom=16'h2FCA;
  11'h128:rom=16'h2704;
  11'h129:rom=16'h2FA9;
  11'h12A:rom=16'hD01;
  11'h12B:rom=16'h1D02;
  11'h12C:rom=16'hF00;
  11'h12D:rom=16'h7102;
  11'h12E:rom=16'hD01;
  11'h12F:rom=16'h2704;
  11'h130:rom=16'h2FCA;
  11'h131:rom=16'h2704;
  11'h132:rom=16'h2FA9;
  11'h133:rom=16'hF00;
  11'h134:rom=16'h2704;
  11'h135:rom=16'h2FA9;
  11'h136:rom=16'hF00;
  11'h137:rom=16'h7103;
  11'h138:rom=16'h2704;
  11'h139:rom=16'h2FA9;
  11'h13A:rom=16'hF00;
  11'h13B:rom=16'h7103;
  11'h13C:rom=16'h2704;
  11'h13D:rom=16'h2FA9;
  11'h13E:rom=16'hF00;
  11'h13F:rom=16'hD01;
  11'h140:rom=16'hD12;
  11'h141:rom=16'h301D;
  11'h142:rom=16'h2123;
  11'h143:rom=16'hD04;
  11'h144:rom=16'hD002;
  11'h145:rom=16'h2120;
  11'h146:rom=16'hD00A;
  11'h147:rom=16'h211E;
  11'h148:rom=16'hD03;
  11'h149:rom=16'h40FF;
  11'h14A:rom=16'h211B;
  11'h14B:rom=16'h3F80;
  11'h14C:rom=16'hE01;
  11'h14D:rom=16'h5008;
  11'h14E:rom=16'h1E01;
  11'h14F:rom=16'h3F90;
  11'h150:rom=16'h2710;
  11'h151:rom=16'h7086;
  11'h152:rom=16'h7101;
  11'h153:rom=16'h2704;
  11'h154:rom=16'h2FCB;
  11'h155:rom=16'h3F80;
  11'h156:rom=16'hE01;
  11'h157:rom=16'h6008;
  11'h158:rom=16'h1E01;
  11'h159:rom=16'h3F90;
  11'h15A:rom=16'hD02;
  11'h15B:rom=16'h8002;
  11'h15C:rom=16'h2710;
  11'h15D:rom=16'hD0D8;
  11'h15E:rom=16'h2903;
  11'h15F:rom=16'h2710;
  11'h160:rom=16'h70B8;
  11'h161:rom=16'h1D02;
  11'h162:rom=16'h7102;
  11'h163:rom=16'h2704;
  11'h164:rom=16'h2FCA;
  11'h165:rom=16'hF00;
  11'h166:rom=16'h27FF;
  11'h167:rom=16'h70FF;
  11'h168:rom=16'h1D0C;
  11'h169:rom=16'h1E06;
  11'h16A:rom=16'hF00;
  11'h16B:rom=16'hC04;
  11'h16C:rom=16'h2704;
  11'h16D:rom=16'h2F53;
  11'h16E:rom=16'h3F90;
  11'h16F:rom=16'hC70;
  11'h170:rom=16'hC61;
  11'h171:rom=16'h2704;
  11'h172:rom=16'hF000;
  11'h173:rom=16'h2702;
  11'h174:rom=16'hC000;
  11'h175:rom=16'h212C;
  11'h176:rom=16'h2704;
  11'h177:rom=16'h2F41;
  11'h178:rom=16'h2701;
  11'h179:rom=16'hC000;
  11'h17A:rom=16'h2127;
  11'h17B:rom=16'h40FF;
  11'h17C:rom=16'hC080;
  11'h17D:rom=16'h2131;
  11'h17E:rom=16'hD0F0;
  11'h17F:rom=16'h210B;
  11'h180:rom=16'hD0E0;
  11'h181:rom=16'h210C;
  11'h182:rom=16'hD0FA;
  11'h183:rom=16'h210D;
  11'h184:rom=16'hD0E1;
  11'h185:rom=16'h211A;
  11'h186:rom=16'hD0AA;
  11'h187:rom=16'h211A;
  11'h188:rom=16'h2704;
  11'h189:rom=16'h2F1A;
  11'h18A:rom=16'h5780;
  11'h18B:rom=16'h2704;
  11'h18C:rom=16'h2F1A;
  11'h18D:rom=16'h5740;
  11'h18E:rom=16'h2704;
  11'h18F:rom=16'h2F1A;
  11'h190:rom=16'h47FD;
  11'h191:rom=16'h7000;
  11'h192:rom=16'hC604;
  11'h193:rom=16'h2902;
  11'h194:rom=16'h5002;
  11'h195:rom=16'hC608;
  11'h196:rom=16'h2902;
  11'h197:rom=16'h5004;
  11'h198:rom=16'hC701;
  11'h199:rom=16'h2102;
  11'h19A:rom=16'h5001;
  11'h19B:rom=16'h2704;
  11'h19C:rom=16'h2F5D;
  11'h19D:rom=16'h2704;
  11'h19E:rom=16'h2F1A;
  11'h19F:rom=16'h2704;
  11'h1A0:rom=16'h2F1A;
  11'h1A1:rom=16'h7500;
  11'h1A2:rom=16'h5702;
  11'h1A3:rom=16'h2704;
  11'h1A4:rom=16'h2F14;
  11'h1A5:rom=16'hC780;
  11'h1A6:rom=16'h2704;
  11'h1A7:rom=16'h290E;
  11'h1A8:rom=16'h6701;
  11'h1A9:rom=16'h5702;
  11'h1AA:rom=16'h2702;
  11'h1AB:rom=16'h2FCD;
  11'h1AC:rom=16'h2704;
  11'h1AD:rom=16'h2F0E;
  11'h1AE:rom=16'hC740;
  11'h1AF:rom=16'h2102;
  11'h1B0:rom=16'h5080;
  11'h1B1:rom=16'h270E;
  11'h1B2:rom=16'h8030;
  11'h1B3:rom=16'h2705;
  11'h1B4:rom=16'h2F5F;
  11'h1B5:rom=16'h3507;
  11'h1B6:rom=16'h2151;
  11'h1B7:rom=16'hC701;
  11'h1B8:rom=16'h210D;
  11'h1B9:rom=16'h2704;
  11'h1BA:rom=16'h2FE7;
  11'h1BB:rom=16'h3005;
  11'h1BC:rom=16'h2109;
  11'h1BD:rom=16'hD1C;
  11'h1BE:rom=16'h3105;
  11'h1BF:rom=16'hC780;
  11'h1C0:rom=16'h2902;
  11'h1C1:rom=16'h3106;
  11'h1C2:rom=16'h1D1C;
  11'h1C3:rom=16'h1E16;
  11'h1C4:rom=16'h2F43;
  11'h1C5:rom=16'h56E0;
  11'h1C6:rom=16'hC580;
  11'h1C7:rom=16'h2903;
  11'h1C8:rom=16'h6640;
  11'h1C9:rom=16'h2F0E;
  11'h1CA:rom=16'hD5FF;
  11'h1CB:rom=16'h21DA;
  11'h1CC:rom=16'h3057;
  11'h1CD:rom=16'h2704;
  11'h1CE:rom=16'h2F7D;
  11'h1CF:rom=16'hC00C;
  11'h1D0:rom=16'h2902;
  11'h1D1:rom=16'h3605;
  11'h1D2:rom=16'hC780;
  11'h1D3:rom=16'h2902;
  11'h1D4:rom=16'h3606;
  11'h1D5:rom=16'h5702;
  11'h1D6:rom=16'h7500;
  11'h1D7:rom=16'hD539;
  11'h1D8:rom=16'h2002;
  11'h1D9:rom=16'h6680;
  11'h1DA:rom=16'hC640;
  11'h1DB:rom=16'h2905;
  11'h1DC:rom=16'hD0B;
  11'h1DD:rom=16'h305D;
  11'h1DE:rom=16'h2902;
  11'h1DF:rom=16'h6620;
  11'h1E0:rom=16'hC780;
  11'h1E1:rom=16'h2108;
  11'h1E2:rom=16'h2704;
  11'h1E3:rom=16'h2F35;
  11'h1E4:rom=16'hC620;
  11'h1E5:rom=16'h2922;
  11'h1E6:rom=16'h5660;
  11'h1E7:rom=16'h7500;
  11'h1E8:rom=16'h1D5B;
  11'h1E9:rom=16'hC640;
  11'h1EA:rom=16'h2902;
  11'h1EB:rom=16'h1D5B;
  11'h1EC:rom=16'h3167;
  11'h1ED:rom=16'h2701;
  11'h1EE:rom=16'hF100;
  11'h1EF:rom=16'h3164;
  11'h1F0:rom=16'h41FF;
  11'h1F1:rom=16'h2705;
  11'h1F2:rom=16'h2F1B;
  11'h1F3:rom=16'h2701;
  11'h1F4:rom=16'hE000;
  11'h1F5:rom=16'h3015;
  11'h1F6:rom=16'hD11;
  11'h1F7:rom=16'hD23;
  11'h1F8:rom=16'h3225;
  11'h1F9:rom=16'h210B;
  11'h1FA:rom=16'h8102;
  11'h1FB:rom=16'h2710;
  11'h1FC:rom=16'hD1D8;
  11'h1FD:rom=16'h2903;
  11'h1FE:rom=16'h2710;
  11'h1FF:rom=16'h71B8;
  11'h200:rom=16'hD22;
  11'h201:rom=16'h321D;
  11'h202:rom=16'h2103;
  11'h203:rom=16'h1D11;
  11'h204:rom=16'h1100;
  11'h205:rom=16'h2704;
  11'h206:rom=16'h2F21;
  11'h207:rom=16'h473F;
  11'h208:rom=16'hC702;
  11'h209:rom=16'h2104;
  11'h20A:rom=16'h70ED;
  11'h20B:rom=16'h2704;
  11'h20C:rom=16'h2F5D;
  11'h20D:rom=16'h1C70;
  11'h20E:rom=16'h1C61;
  11'h20F:rom=16'hF00;
  11'h210:rom=16'hD003;
  11'h211:rom=16'h2909;
  11'h212:rom=16'h3F80;
  11'h213:rom=16'h7001;
  11'h214:rom=16'h2710;
  11'h215:rom=16'h7188;
  11'h216:rom=16'h1100;
  11'h217:rom=16'hE01;
  11'h218:rom=16'h5004;
  11'h219:rom=16'h2F04;
  11'h21A:rom=16'h3F80;
  11'h21B:rom=16'hE01;
  11'h21C:rom=16'h40FB;
  11'h21D:rom=16'h1E01;
  11'h21E:rom=16'h3F90;
  11'h21F:rom=16'hF00;
  11'h220:rom=16'h7101;
  11'h221:rom=16'h301C;
  11'h222:rom=16'h2103;
  11'h223:rom=16'h2701;
  11'h224:rom=16'h6000;
  11'h225:rom=16'h3118;
  11'h226:rom=16'h41FF;
  11'h227:rom=16'h29FA;
  11'h228:rom=16'hF00;
  11'h229:rom=16'h710B;
  11'h22A:rom=16'h1C15;
  11'h22B:rom=16'h7100;
  11'h22C:rom=16'h1C16;
  11'h22D:rom=16'hF00;
  11'h22E:rom=16'h7100;
  11'h22F:rom=16'h1C16;
  11'h230:rom=16'h7180;
  11'h231:rom=16'h1C15;
  11'h232:rom=16'h7101;
  11'h233:rom=16'h1E12;
  11'h234:rom=16'h2701;
  11'h235:rom=16'h5000;
  11'h236:rom=16'h2704;
  11'h237:rom=16'h2F41;
  11'h238:rom=16'h2706;
  11'h239:rom=16'h5000;
  11'h23A:rom=16'h1C04;
  11'h23B:rom=16'h7105;
  11'h23C:rom=16'h1C16;
  11'h23D:rom=16'hF00;
  11'h23E:rom=16'h400F;
  11'h23F:rom=16'h3008;
  11'h240:rom=16'h2704;
  11'h241:rom=16'h8088;
  11'h242:rom=16'h00;
  11'h243:rom=16'hF00;
  11'h244:rom=16'h01;
  11'h245:rom=16'h02;
  11'h246:rom=16'h04;
  11'h247:rom=16'h08;
  11'h248:rom=16'h10;
  11'h249:rom=16'h20;
  11'h24A:rom=16'h40;
  11'h24B:rom=16'h80;
  11'h24C:rom=16'h100;
  11'h24D:rom=16'h200;
  11'h24E:rom=16'h400;
  11'h24F:rom=16'h800;
  11'h250:rom=16'h1000;
  11'h251:rom=16'h2000;
  11'h252:rom=16'h4000;
  11'h253:rom=16'h8000;
  11'h254:rom=16'hE21;
  11'h255:rom=16'hC202;
  11'h256:rom=16'h21FE;
  11'h257:rom=16'hB21;
  11'h258:rom=16'hC001;
  11'h259:rom=16'h2106;
  11'h25A:rom=16'h2701;
  11'h25B:rom=16'hE200;
  11'h25C:rom=16'h30;
  11'h25D:rom=16'h43FF;
  11'h25E:rom=16'h3235;
  11'h25F:rom=16'h1020;
  11'h260:rom=16'hE25;
  11'h261:rom=16'h8001;
  11'h262:rom=16'h9101;
  11'h263:rom=16'h29F1;
  11'h264:rom=16'hF00;
  11'h265:rom=16'h20;
  11'h266:rom=16'hC001;
  11'h267:rom=16'h2103;
  11'h268:rom=16'h2701;
  11'h269:rom=16'hF200;
  11'h26A:rom=16'h1B20;
  11'h26B:rom=16'hE24;
  11'h26C:rom=16'hE21;
  11'h26D:rom=16'hC201;
  11'h26E:rom=16'h29FE;
  11'h26F:rom=16'h8001;
  11'h270:rom=16'h9101;
  11'h271:rom=16'h29F4;
  11'h272:rom=16'hF00;
  11'h273:rom=16'h7001;
  11'h274:rom=16'h2704;
  11'h275:rom=16'h71FA;
  11'h276:rom=16'h120;
  11'h277:rom=16'h325D;
  11'h278:rom=16'h2104;
  11'h279:rom=16'h8102;
  11'h27A:rom=16'h3008;
  11'h27B:rom=16'h29FB;
  11'h27C:rom=16'hF00;
  11'h27D:rom=16'h56;
  11'h27E:rom=16'h50;
  11'h27F:rom=16'h52;
  11'h280:rom=16'h54;
  11'h281:rom=16'h01;
  11'h282:rom=16'h1A;
  11'h283:rom=16'h18;
  11'h284:rom=16'h03;
  11'h285:rom=16'h00;
  11'h286:rom=16'h00;
  11'h287:rom=16'h00;
  11'h288:rom=16'h00;
  11'h289:rom=16'h00;
  11'h28A:rom=16'h00;
  11'h28B:rom=16'h00;
  11'h28C:rom=16'h00;
  11'h28D:rom=16'h3057;
  11'h28E:rom=16'h211E;
  11'h28F:rom=16'hC101;
  11'h290:rom=16'h210D;
  11'h291:rom=16'hD01B;
  11'h292:rom=16'h2010;
  11'h293:rom=16'hC102;
  11'h294:rom=16'h2105;
  11'h295:rom=16'h270F;
  11'h296:rom=16'h8015;
  11'h297:rom=16'h2705;
  11'h298:rom=16'h2F5E;
  11'h299:rom=16'h270F;
  11'h29A:rom=16'h8053;
  11'h29B:rom=16'h2705;
  11'h29C:rom=16'h2F5E;
  11'h29D:rom=16'hD01B;
  11'h29E:rom=16'h2004;
  11'h29F:rom=16'h270F;
  11'h2A0:rom=16'h8091;
  11'h2A1:rom=16'h2F0C;
  11'h2A2:rom=16'h5060;
  11'h2A3:rom=16'hC108;
  11'h2A4:rom=16'h2902;
  11'h2A5:rom=16'h6020;
  11'h2A6:rom=16'hC102;
  11'h2A7:rom=16'h2902;
  11'h2A8:rom=16'h6020;
  11'h2A9:rom=16'hC101;
  11'h2AA:rom=16'h2902;
  11'h2AB:rom=16'h401F;
  11'h2AC:rom=16'hF00;
  11'h2AD:rom=16'h2705;
  11'h2AE:rom=16'h2F5E;
  11'h2AF:rom=16'hC001;
  11'h2B0:rom=16'h2904;
  11'h2B1:rom=16'h00;
  11'h2B2:rom=16'h40FF;
  11'h2B3:rom=16'hF00;
  11'h2B4:rom=16'h00;
  11'h2B5:rom=16'h2701;
  11'h2B6:rom=16'hF000;
  11'h2B7:rom=16'hF00;
  11'h2B8:rom=16'h1F21;
  11'h2B9:rom=16'h2711;
  11'h2BA:rom=16'h7200;
  11'h2BB:rom=16'h1200;
  11'h2BC:rom=16'h1211;
  11'h2BD:rom=16'hF21;
  11'h2BE:rom=16'hF00;
  11'h2BF:rom=16'h27FF;
  11'h2C0:rom=16'h71FF;
  11'h2C1:rom=16'h1D16;
  11'h2C2:rom=16'h2718;
  11'h2C3:rom=16'h7F00;
  11'h2C4:rom=16'h3F02;
  11'h2C5:rom=16'h3F80;
  11'h2C6:rom=16'h1FF1;
  11'h2C7:rom=16'h1F01;
  11'h2C8:rom=16'h1F11;
  11'h2C9:rom=16'h1F21;
  11'h2CA:rom=16'h1F31;
  11'h2CB:rom=16'h1F41;
  11'h2CC:rom=16'h1F51;
  11'h2CD:rom=16'h1F61;
  11'h2CE:rom=16'h1F71;
  11'h2CF:rom=16'h1DF8;
  11'h2D0:rom=16'h2717;
  11'h2D1:rom=16'h7FC0;
  11'h2D2:rom=16'h1F01;
  11'h2D3:rom=16'h7001;
  11'h2D4:rom=16'h2F04;
  11'h2D5:rom=16'h27FF;
  11'h2D6:rom=16'h70FF;
  11'h2D7:rom=16'h2F01;
  11'h2D8:rom=16'h3F80;
  11'h2D9:rom=16'h1D06;
  11'h2DA:rom=16'h1FF1;
  11'h2DB:rom=16'h1F01;
  11'h2DC:rom=16'h1F11;
  11'h2DD:rom=16'h1F21;
  11'h2DE:rom=16'h1F31;
  11'h2DF:rom=16'h1F41;
  11'h2E0:rom=16'h1F51;
  11'h2E1:rom=16'h1F61;
  11'h2E2:rom=16'h1F71;
  11'h2E3:rom=16'h1DF7;
  11'h2E4:rom=16'hDF8;
  11'h2E5:rom=16'hF71;
  11'h2E6:rom=16'hF61;
  11'h2E7:rom=16'hF51;
  11'h2E8:rom=16'hF41;
  11'h2E9:rom=16'hF31;
  11'h2EA:rom=16'hF21;
  11'h2EB:rom=16'hF11;
  11'h2EC:rom=16'hF01;
  11'h2ED:rom=16'hFF1;
  11'h2EE:rom=16'hF90;
  11'h2EF:rom=16'h3F80;
  11'h2F0:rom=16'hD06;
  11'h2F1:rom=16'hD000;
  11'h2F2:rom=16'h2902;
  11'h2F3:rom=16'hF90;
  11'h2F4:rom=16'h7000;
  11'h2F5:rom=16'h1D06;
  11'h2F6:rom=16'h1FF1;
  11'h2F7:rom=16'h1F01;
  11'h2F8:rom=16'h2F07;
  11'h2F9:rom=16'h1F01;
  11'h2FA:rom=16'hD06;
  11'h2FB:rom=16'h9001;
  11'h2FC:rom=16'h2313;
  11'h2FD:rom=16'h1D06;
  11'h2FE:rom=16'h2911;
  11'h2FF:rom=16'h1F11;
  11'h300:rom=16'h1F21;
  11'h301:rom=16'h1F31;
  11'h302:rom=16'h1F41;
  11'h303:rom=16'h1F51;
  11'h304:rom=16'h1F61;
  11'h305:rom=16'h1F71;
  11'h306:rom=16'h1DF8;
  11'h307:rom=16'hDF7;
  11'h308:rom=16'hF71;
  11'h309:rom=16'hF61;
  11'h30A:rom=16'hF51;
  11'h30B:rom=16'hF41;
  11'h30C:rom=16'hF31;
  11'h30D:rom=16'hF21;
  11'h30E:rom=16'hF11;
  11'h30F:rom=16'hF01;
  11'h310:rom=16'hFF1;
  11'h311:rom=16'hF90;
  11'h312:rom=16'h1FF1;
  11'h313:rom=16'h1F01;
  11'h314:rom=16'hB08;
  11'h315:rom=16'h40FF;
  11'h316:rom=16'h1B08;
  11'h317:rom=16'h7001;
  11'h318:rom=16'h2705;
  11'h319:rom=16'h2FDF;
  11'h31A:rom=16'hF01;
  11'h31B:rom=16'hFF1;
  11'h31C:rom=16'hF90;
  11'h31D:rom=16'h7000;
  11'h31E:rom=16'h1E03;
  11'h31F:rom=16'hE07;
  11'h320:rom=16'h270A;
  11'h321:rom=16'h2FE3;
  11'h322:rom=16'h2780;
  11'h323:rom=16'h7000;
  11'h324:rom=16'h1B08;
  11'h325:rom=16'h7600;
  11'h326:rom=16'h7700;
  11'h327:rom=16'hE13;
  11'h328:rom=16'h41FE;
  11'h329:rom=16'h1E13;
  11'h32A:rom=16'hB08;
  11'h32B:rom=16'h300C;
  11'h32C:rom=16'h2B0A;
  11'h32D:rom=16'h2708;
  11'h32E:rom=16'h2FCF;
  11'h32F:rom=16'h7010;
  11'h330:rom=16'h2705;
  11'h331:rom=16'h2FB1;
  11'h332:rom=16'h2FF8;
  11'h333:rom=16'h70A0;
  11'h334:rom=16'h9001;
  11'h335:rom=16'h29FF;
  11'h336:rom=16'h3707;
  11'h337:rom=16'h2780;
  11'h338:rom=16'h7000;
  11'h339:rom=16'h1B08;
  11'h33A:rom=16'hC780;
  11'h33B:rom=16'h2108;
  11'h33C:rom=16'hC740;
  11'h33D:rom=16'h216D;
  11'h33E:rom=16'hD7F0;
  11'h33F:rom=16'h2708;
  11'h340:rom=16'h20EE;
  11'h341:rom=16'h2708;
  11'h342:rom=16'h2FFC;
  11'h343:rom=16'hE03;
  11'h344:rom=16'h4080;
  11'h345:rom=16'h5001;
  11'h346:rom=16'h1E03;
  11'h347:rom=16'hE07;
  11'h348:rom=16'h2708;
  11'h349:rom=16'h2FCF;
  11'h34A:rom=16'h46F7;
  11'h34B:rom=16'hC708;
  11'h34C:rom=16'h2102;
  11'h34D:rom=16'h5608;
  11'h34E:rom=16'h70BB;
  11'h34F:rom=16'h2705;
  11'h350:rom=16'h2FB1;
  11'h351:rom=16'hC740;
  11'h352:rom=16'h2912;
  11'h353:rom=16'hC720;
  11'h354:rom=16'h2914;
  11'h355:rom=16'hC710;
  11'h356:rom=16'h2906;
  11'h357:rom=16'h71FF;
  11'h358:rom=16'h1B19;
  11'h359:rom=16'h7100;
  11'h35A:rom=16'h1B1B;
  11'h35B:rom=16'h5710;
  11'h35C:rom=16'h5610;
  11'h35D:rom=16'hB0B;
  11'h35E:rom=16'hB19;
  11'h35F:rom=16'h301D;
  11'h360:rom=16'h212D;
  11'h361:rom=16'h2802;
  11'h362:rom=16'h6610;
  11'h363:rom=16'h2F07;
  11'h364:rom=16'h5610;
  11'h365:rom=16'hC720;
  11'h366:rom=16'h2102;
  11'h367:rom=16'h6610;
  11'h368:rom=16'hC710;
  11'h369:rom=16'h2107;
  11'h36A:rom=16'hB09;
  11'h36B:rom=16'h8001;
  11'h36C:rom=16'hC610;
  11'h36D:rom=16'h2902;
  11'h36E:rom=16'h9002;
  11'h36F:rom=16'h1B09;
  11'h370:rom=16'h2708;
  11'h371:rom=16'h2FCF;
  11'h372:rom=16'hC610;
  11'h373:rom=16'h2907;
  11'h374:rom=16'hE03;
  11'h375:rom=16'hC004;
  11'h376:rom=16'h2104;
  11'h377:rom=16'h7000;
  11'h378:rom=16'h1B09;
  11'h379:rom=16'h2F14;
  11'h37A:rom=16'h2709;
  11'h37B:rom=16'h2F31;
  11'h37C:rom=16'h2701;
  11'h37D:rom=16'h7077;
  11'h37E:rom=16'hC703;
  11'h37F:rom=16'h210A;
  11'h380:rom=16'h3008;
  11'h381:rom=16'hC702;
  11'h382:rom=16'h2107;
  11'h383:rom=16'h2704;
  11'h384:rom=16'h70E2;
  11'h385:rom=16'hC701;
  11'h386:rom=16'h2103;
  11'h387:rom=16'h2707;
  11'h388:rom=16'h7053;
  11'h389:rom=16'h2705;
  11'h38A:rom=16'h2FB1;
  11'h38B:rom=16'hC7E0;
  11'h38C:rom=16'h21D0;
  11'h38D:rom=16'hC704;
  11'h38E:rom=16'h210C;
  11'h38F:rom=16'h2707;
  11'h390:rom=16'h2F37;
  11'h391:rom=16'h7000;
  11'h392:rom=16'h1A00;
  11'h393:rom=16'h2708;
  11'h394:rom=16'h2F81;
  11'h395:rom=16'h2707;
  11'h396:rom=16'h3034;
  11'h397:rom=16'hE13;
  11'h398:rom=16'h41F7;
  11'h399:rom=16'h1E13;
  11'h39A:rom=16'h2F8D;
  11'h39B:rom=16'hC704;
  11'h39C:rom=16'h2105;
  11'h39D:rom=16'h2703;
  11'h39E:rom=16'h70A9;
  11'h39F:rom=16'h2705;
  11'h3A0:rom=16'h2FB1;
  11'h3A1:rom=16'h5608;
  11'h3A2:rom=16'hF00;
  11'h3A3:rom=16'h2706;
  11'h3A4:rom=16'h2F4E;
  11'h3A5:rom=16'hE13;
  11'h3A6:rom=16'h5140;
  11'h3A7:rom=16'h1E13;
  11'h3A8:rom=16'h2706;
  11'h3A9:rom=16'h2F4E;
  11'h3AA:rom=16'hE03;
  11'h3AB:rom=16'h4080;
  11'h3AC:rom=16'h5001;
  11'h3AD:rom=16'h1E03;
  11'h3AE:rom=16'h2708;
  11'h3AF:rom=16'h2FCF;
  11'h3B0:rom=16'h7010;
  11'h3B1:rom=16'h2705;
  11'h3B2:rom=16'h2FB1;
  11'h3B3:rom=16'hE03;
  11'h3B4:rom=16'hC080;
  11'h3B5:rom=16'h29EE;
  11'h3B6:rom=16'h5608;
  11'h3B7:rom=16'hC704;
  11'h3B8:rom=16'h2105;
  11'h3B9:rom=16'h2703;
  11'h3BA:rom=16'h70A9;
  11'h3BB:rom=16'h2705;
  11'h3BC:rom=16'h2FB1;
  11'h3BD:rom=16'h2708;
  11'h3BE:rom=16'h2F6D;
  11'h3BF:rom=16'h46FE;
  11'h3C0:rom=16'hB09;
  11'h3C1:rom=16'hD02C;
  11'h3C2:rom=16'h2002;
  11'h3C3:rom=16'h5601;
  11'h3C4:rom=16'hC720;
  11'h3C5:rom=16'h2104;
  11'h3C6:rom=16'hE03;
  11'h3C7:rom=16'h2702;
  11'h3C8:rom=16'hC000;
  11'h3C9:rom=16'h7000;
  11'h3CA:rom=16'h1A00;
  11'h3CB:rom=16'h2708;
  11'h3CC:rom=16'h2F81;
  11'h3CD:rom=16'h2042;
  11'h3CE:rom=16'hB08;
  11'h3CF:rom=16'h300C;
  11'h3D0:rom=16'h2706;
  11'h3D1:rom=16'h2B6C;
  11'h3D2:rom=16'hC702;
  11'h3D3:rom=16'h2107;
  11'h3D4:rom=16'hA05;
  11'h3D5:rom=16'hC708;
  11'h3D6:rom=16'h2102;
  11'h3D7:rom=16'h6001;
  11'h3D8:rom=16'hC001;
  11'h3D9:rom=16'h29F2;
  11'h3DA:rom=16'hA06;
  11'h3DB:rom=16'hB1A;
  11'h3DC:rom=16'h301D;
  11'h3DD:rom=16'h29EE;
  11'h3DE:rom=16'hA08;
  11'h3DF:rom=16'hC008;
  11'h3E0:rom=16'h2105;
  11'h3E1:rom=16'hE03;
  11'h3E2:rom=16'h5008;
  11'h3E3:rom=16'h1E03;
  11'h3E4:rom=16'h2FE7;
  11'h3E5:rom=16'hE03;
  11'h3E6:rom=16'h40F7;
  11'h3E7:rom=16'h1E03;
  11'h3E8:rom=16'hC720;
  11'h3E9:rom=16'h2928;
  11'h3EA:rom=16'hA1A;
  11'h3EB:rom=16'hA2B;
  11'h3EC:rom=16'h2751;
  11'h3ED:rom=16'h5200;
  11'h3EE:rom=16'hA31;
  11'h3EF:rom=16'h7002;
  11'h3F0:rom=16'h2705;
  11'h3F1:rom=16'h2FB1;
  11'h3F2:rom=16'h3F80;
  11'h3F3:rom=16'h1E18;
  11'h3F4:rom=16'h1E29;
  11'h3F5:rom=16'h8101;
  11'h3F6:rom=16'hA200;
  11'h3F7:rom=16'hE00;
  11'h3F8:rom=16'h2702;
  11'h3F9:rom=16'hC000;
  11'h3FA:rom=16'h29FD;
  11'h3FB:rom=16'hE00;
  11'h3FC:rom=16'h40FF;
  11'h3FD:rom=16'h1B0B;
  11'h3FE:rom=16'h7000;
  11'h3FF:rom=16'h1E09;
  11'h400:rom=16'h3F90;
  11'h401:rom=16'hE06;
  11'h402:rom=16'h9301;
  11'h403:rom=16'h29EC;
  11'h404:rom=16'h7004;
  11'h405:rom=16'h2705;
  11'h406:rom=16'h2FB1;
  11'h407:rom=16'hC710;
  11'h408:rom=16'h2706;
  11'h409:rom=16'h214E;
  11'h40A:rom=16'hB0A;
  11'h40B:rom=16'h8001;
  11'h40C:rom=16'h40FF;
  11'h40D:rom=16'h1B0A;
  11'h40E:rom=16'h2FBB;
  11'h40F:rom=16'h2706;
  11'h410:rom=16'h2F4E;
  11'h411:rom=16'hE06;
  11'h412:rom=16'hC701;
  11'h413:rom=16'h7002;
  11'h414:rom=16'h2705;
  11'h415:rom=16'h2FB1;
  11'h416:rom=16'h3F80;
  11'h417:rom=16'hB0B;
  11'h418:rom=16'h1E00;
  11'h419:rom=16'h1F11;
  11'h41A:rom=16'hA0A;
  11'h41B:rom=16'h1E08;
  11'h41C:rom=16'hA1B;
  11'h41D:rom=16'h2791;
  11'h41E:rom=16'h5100;
  11'h41F:rom=16'h1E19;
  11'h420:rom=16'h8001;
  11'h421:rom=16'hA100;
  11'h422:rom=16'h1A1B;
  11'h423:rom=16'h1A0A;
  11'h424:rom=16'hF11;
  11'h425:rom=16'hE00;
  11'h426:rom=16'h2702;
  11'h427:rom=16'hC000;
  11'h428:rom=16'h29FD;
  11'h429:rom=16'h7000;
  11'h42A:rom=16'h1E09;
  11'h42B:rom=16'h3F90;
  11'h42C:rom=16'hA01;
  11'h42D:rom=16'h9001;
  11'h42E:rom=16'h1A01;
  11'h42F:rom=16'h2103;
  11'h430:rom=16'hE06;
  11'h431:rom=16'h2FE2;
  11'h432:rom=16'h7004;
  11'h433:rom=16'h2705;
  11'h434:rom=16'h2FB1;
  11'h435:rom=16'h2FD2;
  11'h436:rom=16'hF00;
  11'h437:rom=16'hE03;
  11'h438:rom=16'h2701;
  11'h439:rom=16'hC000;
  11'h43A:rom=16'h2102;
  11'h43B:rom=16'hF00;
  11'h43C:rom=16'h7002;
  11'h43D:rom=16'h2705;
  11'h43E:rom=16'h2FB1;
  11'h43F:rom=16'h2FF7;
  11'h440:rom=16'hA00;
  11'h441:rom=16'hD005;
  11'h442:rom=16'h2820;
  11'h443:rom=16'h2709;
  11'h444:rom=16'h2F8B;
  11'h445:rom=16'h201C;
  11'h446:rom=16'hA17;
  11'h447:rom=16'h7080;
  11'h448:rom=16'h9101;
  11'h449:rom=16'h2008;
  11'h44A:rom=16'h3008;
  11'h44B:rom=16'h9101;
  11'h44C:rom=16'h2005;
  11'h44D:rom=16'h3008;
  11'h44E:rom=16'h9101;
  11'h44F:rom=16'h2002;
  11'h450:rom=16'h3008;
  11'h451:rom=16'h1A01;
  11'h452:rom=16'h2708;
  11'h453:rom=16'h2FCF;
  11'h454:rom=16'hB09;
  11'h455:rom=16'hA14;
  11'h456:rom=16'h301D;
  11'h457:rom=16'h2108;
  11'h458:rom=16'hA01;
  11'h459:rom=16'h804E;
  11'h45A:rom=16'h2701;
  11'h45B:rom=16'hF000;
  11'h45C:rom=16'h2705;
  11'h45D:rom=16'h2FB1;
  11'h45E:rom=16'h2FE2;
  11'h45F:rom=16'h3F20;
  11'h460:rom=16'hF00;
  11'h461:rom=16'h2FDF;
  11'h462:rom=16'hE13;
  11'h463:rom=16'h5110;
  11'h464:rom=16'h1E13;
  11'h465:rom=16'h3F30;
  11'h466:rom=16'hF00;
  11'h467:rom=16'h2709;
  11'h468:rom=16'h2F4B;
  11'h469:rom=16'h70C8;
  11'h46A:rom=16'hC780;
  11'h46B:rom=16'h2902;
  11'h46C:rom=16'h70C6;
  11'h46D:rom=16'h3F80;
  11'h46E:rom=16'hA18;
  11'h46F:rom=16'h3104;
  11'h470:rom=16'hE23;
  11'h471:rom=16'h3205;
  11'h472:rom=16'h3206;
  11'h473:rom=16'h3125;
  11'h474:rom=16'h1E13;
  11'h475:rom=16'h3F90;
  11'h476:rom=16'hF00;
  11'h477:rom=16'h27FF;
  11'h478:rom=16'h70F0;
  11'h479:rom=16'h1E07;
  11'h47A:rom=16'h3F80;
  11'h47B:rom=16'h2FFC;
  11'h47C:rom=16'h2706;
  11'h47D:rom=16'h2F4E;
  11'h47E:rom=16'h2706;
  11'h47F:rom=16'h2F4E;
  11'h480:rom=16'hB0C;
  11'h481:rom=16'hA18;
  11'h482:rom=16'hC080;
  11'h483:rom=16'h210E;
  11'h484:rom=16'hC002;
  11'h485:rom=16'h290C;
  11'h486:rom=16'h4001;
  11'h487:rom=16'h3107;
  11'h488:rom=16'h8101;
  11'h489:rom=16'h1E14;
  11'h48A:rom=16'hE006;
  11'h48B:rom=16'h2710;
  11'h48C:rom=16'h80F4;
  11'h48D:rom=16'h417F;
  11'h48E:rom=16'h1A0D;
  11'h48F:rom=16'h1A18;
  11'h490:rom=16'hF00;
  11'h491:rom=16'h7000;
  11'h492:rom=16'h1E04;
  11'h493:rom=16'h2710;
  11'h494:rom=16'h70F4;
  11'h495:rom=16'h5180;
  11'h496:rom=16'h21FB;
  11'h497:rom=16'h2FF7;
  11'h498:rom=16'h7000;
  11'h499:rom=16'h71A0;
  11'h49A:rom=16'h2705;
  11'h49B:rom=16'h2F71;
  11'h49C:rom=16'h2709;
  11'h49D:rom=16'h2F01;
  11'h49E:rom=16'h10;
  11'h49F:rom=16'h8101;
  11'h4A0:rom=16'hC610;
  11'h4A1:rom=16'h2902;
  11'h4A2:rom=16'h9102;
  11'h4A3:rom=16'h1010;
  11'h4A4:rom=16'h2F04;
  11'h4A5:rom=16'h2709;
  11'h4A6:rom=16'h2F01;
  11'h4A7:rom=16'h10;
  11'h4A8:rom=16'hD101;
  11'h4A9:rom=16'h2807;
  11'h4AA:rom=16'h7100;
  11'h4AB:rom=16'h1010;
  11'h4AC:rom=16'hA08;
  11'h4AD:rom=16'h5004;
  11'h4AE:rom=16'h1A08;
  11'h4AF:rom=16'hF00;
  11'h4B0:rom=16'hD12B;
  11'h4B1:rom=16'h2003;
  11'h4B2:rom=16'h712B;
  11'h4B3:rom=16'h1010;
  11'h4B4:rom=16'hA08;
  11'h4B5:rom=16'h40FB;
  11'h4B6:rom=16'h1A08;
  11'h4B7:rom=16'hF00;
  11'h4B8:rom=16'h2709;
  11'h4B9:rom=16'h2F01;
  11'h4BA:rom=16'h11;
  11'h4BB:rom=16'h22;
  11'h4BC:rom=16'h1A1A;
  11'h4BD:rom=16'h1A2B;
  11'h4BE:rom=16'h00;
  11'h4BF:rom=16'h3008;
  11'h4C0:rom=16'hB1C;
  11'h4C1:rom=16'hC110;
  11'h4C2:rom=16'h2102;
  11'h4C3:rom=16'h5001;
  11'h4C4:rom=16'hF00;
  11'h4C5:rom=16'h2709;
  11'h4C6:rom=16'h2F71;
  11'h4C7:rom=16'h270A;
  11'h4C8:rom=16'h2F5D;
  11'h4C9:rom=16'h282A;
  11'h4CA:rom=16'h2709;
  11'h4CB:rom=16'h2F71;
  11'h4CC:rom=16'h3107;
  11'h4CD:rom=16'h2780;
  11'h4CE:rom=16'hF100;
  11'h4CF:rom=16'h1A14;
  11'h4D0:rom=16'h3107;
  11'h4D1:rom=16'h4101;
  11'h4D2:rom=16'h1A15;
  11'h4D3:rom=16'hA29;
  11'h4D4:rom=16'h8201;
  11'h4D5:rom=16'hD210;
  11'h4D6:rom=16'h2005;
  11'h4D7:rom=16'hA20;
  11'h4D8:rom=16'h8201;
  11'h4D9:rom=16'h1A20;
  11'h4DA:rom=16'h7200;
  11'h4DB:rom=16'h1A29;
  11'h4DC:rom=16'h8201;
  11'h4DD:rom=16'h1A26;
  11'h4DE:rom=16'h9201;
  11'h4DF:rom=16'hE010;
  11'h4E0:rom=16'h3028;
  11'h4E1:rom=16'h3107;
  11'h4E2:rom=16'h2701;
  11'h4E3:rom=16'hE000;
  11'h4E4:rom=16'h2701;
  11'h4E5:rom=16'hF100;
  11'h4E6:rom=16'hA2A;
  11'h4E7:rom=16'h3028;
  11'h4E8:rom=16'hA2B;
  11'h4E9:rom=16'h312A;
  11'h4EA:rom=16'h1A0A;
  11'h4EB:rom=16'h1A1B;
  11'h4EC:rom=16'hA08;
  11'h4ED:rom=16'h40C7;
  11'h4EE:rom=16'h1A08;
  11'h4EF:rom=16'h7001;
  11'h4F0:rom=16'h1A07;
  11'h4F1:rom=16'h3F20;
  11'h4F2:rom=16'hF00;
  11'h4F3:rom=16'h2709;
  11'h4F4:rom=16'h2F71;
  11'h4F5:rom=16'hE004;
  11'h4F6:rom=16'h8020;
  11'h4F7:rom=16'hA2A;
  11'h4F8:rom=16'hA1B;
  11'h4F9:rom=16'h3028;
  11'h4FA:rom=16'hA100;
  11'h4FB:rom=16'h270A;
  11'h4FC:rom=16'h2FCD;
  11'h4FD:rom=16'h3327;
  11'h4FE:rom=16'h270A;
  11'h4FF:rom=16'h2FCD;
  11'h500:rom=16'hA0A;
  11'h501:rom=16'hA1B;
  11'h502:rom=16'h3038;
  11'h503:rom=16'h312A;
  11'h504:rom=16'h8004;
  11'h505:rom=16'hA100;
  11'h506:rom=16'h270A;
  11'h507:rom=16'h2FCD;
  11'h508:rom=16'h9006;
  11'h509:rom=16'hB100;
  11'h50A:rom=16'hA39;
  11'h50B:rom=16'h8301;
  11'h50C:rom=16'h332D;
  11'h50D:rom=16'h2005;
  11'h50E:rom=16'hA30;
  11'h50F:rom=16'h8301;
  11'h510:rom=16'h1A30;
  11'h511:rom=16'h7300;
  11'h512:rom=16'h1A39;
  11'h513:rom=16'h9301;
  11'h514:rom=16'h2008;
  11'h515:rom=16'h800E;
  11'h516:rom=16'hA100;
  11'h517:rom=16'h270A;
  11'h518:rom=16'h2FCD;
  11'h519:rom=16'h3028;
  11'h51A:rom=16'hA100;
  11'h51B:rom=16'h2FF8;
  11'h51C:rom=16'h270A;
  11'h51D:rom=16'h2FAD;
  11'h51E:rom=16'h1A24;
  11'h51F:rom=16'h270A;
  11'h520:rom=16'h2FAD;
  11'h521:rom=16'h1A25;
  11'h522:rom=16'h270A;
  11'h523:rom=16'h2FAD;
  11'h524:rom=16'h1A26;
  11'h525:rom=16'h270A;
  11'h526:rom=16'h2FAD;
  11'h527:rom=16'h1A27;
  11'h528:rom=16'h800C;
  11'h529:rom=16'hA100;
  11'h52A:rom=16'h1A0A;
  11'h52B:rom=16'h1A1B;
  11'h52C:rom=16'hF00;
  11'h52D:rom=16'hF00;
  11'h52E:rom=16'h270A;
  11'h52F:rom=16'h2F5B;
  11'h530:rom=16'hA0A;
  11'h531:rom=16'hA1B;
  11'h532:rom=16'h721A;
  11'h533:rom=16'h3028;
  11'h534:rom=16'hA100;
  11'h535:rom=16'h270A;
  11'h536:rom=16'h2FAD;
  11'h537:rom=16'hD200;
  11'h538:rom=16'h2104;
  11'h539:rom=16'hA38;
  11'h53A:rom=16'h5340;
  11'h53B:rom=16'h1A38;
  11'h53C:rom=16'h270A;
  11'h53D:rom=16'h2FAD;
  11'h53E:rom=16'hD200;
  11'h53F:rom=16'h2106;
  11'h540:rom=16'hD210;
  11'h541:rom=16'h2104;
  11'h542:rom=16'hD220;
  11'h543:rom=16'h2102;
  11'h544:rom=16'h2F0E;
  11'h545:rom=16'h8004;
  11'h546:rom=16'hA100;
  11'h547:rom=16'h270A;
  11'h548:rom=16'h2FCD;
  11'h549:rom=16'h2702;
  11'h54A:rom=16'hD2B0;
  11'h54B:rom=16'h2907;
  11'h54C:rom=16'h270A;
  11'h54D:rom=16'h2FCD;
  11'h54E:rom=16'hD200;
  11'h54F:rom=16'h2903;
  11'h550:rom=16'h3F20;
  11'h551:rom=16'hF00;
  11'h552:rom=16'h270A;
  11'h553:rom=16'h2F5B;
  11'h554:rom=16'h3F30;
  11'h555:rom=16'hF00;
  11'h556:rom=16'h3F80;
  11'h557:rom=16'h1E08;
  11'h558:rom=16'h2751;
  11'h559:rom=16'h5100;
  11'h55A:rom=16'h1E19;
  11'h55B:rom=16'h8001;
  11'h55C:rom=16'hA100;
  11'h55D:rom=16'hE20;
  11'h55E:rom=16'h2702;
  11'h55F:rom=16'hC200;
  11'h560:rom=16'h29FD;
  11'h561:rom=16'hE20;
  11'h562:rom=16'h42FF;
  11'h563:rom=16'h1E29;
  11'h564:rom=16'h3F90;
  11'h565:rom=16'hF00;
  11'h566:rom=16'h1F31;
  11'h567:rom=16'h270A;
  11'h568:rom=16'h2FAD;
  11'h569:rom=16'h3327;
  11'h56A:rom=16'h270A;
  11'h56B:rom=16'h2FAD;
  11'h56C:rom=16'h2701;
  11'h56D:rom=16'hE200;
  11'h56E:rom=16'h3235;
  11'h56F:rom=16'hF31;
  11'h570:rom=16'hF00;
  11'h571:rom=16'h7000;
  11'h572:rom=16'h1B09;
  11'h573:rom=16'h7001;
  11'h574:rom=16'h1B0A;
  11'h575:rom=16'h7010;
  11'h576:rom=16'h1B0B;
  11'h577:rom=16'h7080;
  11'h578:rom=16'h1B0C;
  11'h579:rom=16'h7000;
  11'h57A:rom=16'h1A08;
  11'h57B:rom=16'h2710;
  11'h57C:rom=16'h72F4;
  11'h57D:rom=16'h7000;
  11'h57E:rom=16'h7101;
  11'h57F:rom=16'h270B;
  11'h580:rom=16'h2F0D;
  11'h581:rom=16'h2710;
  11'h582:rom=16'h72FA;
  11'h583:rom=16'h2780;
  11'h584:rom=16'h7000;
  11'h585:rom=16'h7107;
  11'h586:rom=16'h1201;
  11'h587:rom=16'h1212;
  11'h588:rom=16'h7000;
  11'h589:rom=16'h1200;
  11'h58A:rom=16'hF00;
  11'h58B:rom=16'h1FF1;
  11'h58C:rom=16'h1F01;
  11'h58D:rom=16'h1F11;
  11'h58E:rom=16'h1F71;
  11'h58F:rom=16'hB03;
  11'h590:rom=16'h3005;
  11'h591:rom=16'h2308;
  11'h592:rom=16'h2780;
  11'h593:rom=16'h7100;
  11'h594:rom=16'h1B13;
  11'h595:rom=16'h2711;
  11'h596:rom=16'h772E;
  11'h597:rom=16'h710;
  11'h598:rom=16'h3F13;
  11'h599:rom=16'hE00;
  11'h59A:rom=16'h2704;
  11'h59B:rom=16'hC000;
  11'h59C:rom=16'h2103;
  11'h59D:rom=16'h270D;
  11'h59E:rom=16'h2F29;
  11'h59F:rom=16'hF71;
  11'h5A0:rom=16'hF11;
  11'h5A1:rom=16'hF01;
  11'h5A2:rom=16'hFF1;
  11'h5A3:rom=16'hF90;
  11'h5A4:rom=16'h716;
  11'h5A5:rom=16'h41FE;
  11'h5A6:rom=16'h1716;
  11'h5A7:rom=16'h714;
  11'h5A8:rom=16'h41BF;
  11'h5A9:rom=16'h1714;
  11'h5AA:rom=16'hF00;
  11'h5AB:rom=16'h714;
  11'h5AC:rom=16'h5140;
  11'h5AD:rom=16'h1714;
  11'h5AE:rom=16'h706;
  11'h5AF:rom=16'h714;
  11'h5B0:rom=16'h3015;
  11'h5B1:rom=16'h1E0A;
  11'h5B2:rom=16'hF00;
  11'h5B3:rom=16'h716;
  11'h5B4:rom=16'h5101;
  11'h5B5:rom=16'h2FF1;
  11'h5B6:rom=16'h270B;
  11'h5B7:rom=16'h7174;
  11'h5B8:rom=16'h1710;
  11'h5B9:rom=16'h2FED;
  11'h5BA:rom=16'h2F61;
  11'h5BB:rom=16'h2711;
  11'h5BC:rom=16'h711A;
  11'h5BD:rom=16'h708;
  11'h5BE:rom=16'h1102;
  11'h5BF:rom=16'h709;
  11'h5C0:rom=16'h1103;
  11'h5C1:rom=16'h1F21;
  11'h5C2:rom=16'h1F31;
  11'h5C3:rom=16'h2711;
  11'h5C4:rom=16'h711A;
  11'h5C5:rom=16'h2711;
  11'h5C6:rom=16'h721C;
  11'h5C7:rom=16'h3317;
  11'h5C8:rom=16'h701;
  11'h5C9:rom=16'hC004;
  11'h5CA:rom=16'h2903;
  11'h5CB:rom=16'h8102;
  11'h5CC:rom=16'h9202;
  11'h5CD:rom=16'h1318;
  11'h5CE:rom=16'h1329;
  11'h5CF:rom=16'h1F21;
  11'h5D0:rom=16'h3217;
  11'h5D1:rom=16'h270D;
  11'h5D2:rom=16'h2FD9;
  11'h5D3:rom=16'h2740;
  11'h5D4:rom=16'h5000;
  11'h5D5:rom=16'h1204;
  11'h5D6:rom=16'hF21;
  11'h5D7:rom=16'h270D;
  11'h5D8:rom=16'h2FD9;
  11'h5D9:rom=16'h2780;
  11'h5DA:rom=16'h5000;
  11'h5DB:rom=16'h1204;
  11'h5DC:rom=16'hF31;
  11'h5DD:rom=16'hF21;
  11'h5DE:rom=16'h2711;
  11'h5DF:rom=16'h711A;
  11'h5E0:rom=16'h70A;
  11'h5E1:rom=16'h3005;
  11'h5E2:rom=16'h2902;
  11'h5E3:rom=16'h9001;
  11'h5E4:rom=16'h1101;
  11'h5E5:rom=16'h2FBF;
  11'h5E6:rom=16'h1707;
  11'h5E7:rom=16'hD0D4;
  11'h5E8:rom=16'h28BC;
  11'h5E9:rom=16'h2780;
  11'h5EA:rom=16'hF000;
  11'h5EB:rom=16'h403E;
  11'h5EC:rom=16'h270B;
  11'h5ED:rom=16'h80E0;
  11'h5EE:rom=16'h00;
  11'h5EF:rom=16'h3F02;
  11'h5F0:rom=16'hB48;
  11'h5F1:rom=16'hB56;
  11'h5F2:rom=16'hB48;
  11'h5F3:rom=16'hB48;
  11'h5F4:rom=16'hB48;
  11'h5F5:rom=16'hB48;
  11'h5F6:rom=16'hB48;
  11'h5F7:rom=16'hB48;
  11'h5F8:rom=16'hB48;
  11'h5F9:rom=16'hB48;
  11'h5FA:rom=16'hB48;
  11'h5FB:rom=16'hB48;
  11'h5FC:rom=16'hB66;
  11'h5FD:rom=16'hB48;
  11'h5FE:rom=16'hB6C;
  11'h5FF:rom=16'hB48;
  11'h600:rom=16'hB48;
  11'h601:rom=16'hB48;
  11'h602:rom=16'hB48;
  11'h603:rom=16'hB76;
  11'h604:rom=16'hB82;
  11'h605:rom=16'hC087;
  11'h606:rom=16'h211E;
  11'h607:rom=16'hC083;
  11'h608:rom=16'h210E;
  11'h609:rom=16'hC080;
  11'h60A:rom=16'h2115;
  11'h60B:rom=16'hC003;
  11'h60C:rom=16'h211C;
  11'h60D:rom=16'hC002;
  11'h60E:rom=16'h2123;
  11'h60F:rom=16'hC001;
  11'h610:rom=16'h270B;
  11'h611:rom=16'h29CC;
  11'h612:rom=16'h270C;
  11'h613:rom=16'h71B6;
  11'h614:rom=16'h1706;
  11'h615:rom=16'hF00;
  11'h616:rom=16'h1702;
  11'h617:rom=16'h270C;
  11'h618:rom=16'h71B2;
  11'h619:rom=16'hC040;
  11'h61A:rom=16'h2903;
  11'h61B:rom=16'h270C;
  11'h61C:rom=16'h710A;
  11'h61D:rom=16'h1710;
  11'h61E:rom=16'hF00;
  11'h61F:rom=16'h1701;
  11'h620:rom=16'h270C;
  11'h621:rom=16'h716C;
  11'h622:rom=16'hC078;
  11'h623:rom=16'h2FF7;
  11'h624:rom=16'h1703;
  11'h625:rom=16'h270C;
  11'h626:rom=16'h71B6;
  11'h627:rom=16'h2FF2;
  11'h628:rom=16'h1704;
  11'h629:rom=16'hC040;
  11'h62A:rom=16'h2103;
  11'h62B:rom=16'h270B;
  11'h62C:rom=16'h2F5D;
  11'h62D:rom=16'h270C;
  11'h62E:rom=16'h71BA;
  11'h62F:rom=16'hC018;
  11'h630:rom=16'h2FEA;
  11'h631:rom=16'h1705;
  11'h632:rom=16'h270C;
  11'h633:rom=16'h71CC;
  11'h634:rom=16'hC01C;
  11'h635:rom=16'h2FE5;
  11'h636:rom=16'h3107;
  11'h637:rom=16'h701;
  11'h638:rom=16'hC008;
  11'h639:rom=16'h2108;
  11'h63A:rom=16'h6008;
  11'h63B:rom=16'h728;
  11'h63C:rom=16'h27FF;
  11'h63D:rom=16'h4200;
  11'h63E:rom=16'h3215;
  11'h63F:rom=16'h1728;
  11'h640:rom=16'h2FDF;
  11'h641:rom=16'hC010;
  11'h642:rom=16'h2107;
  11'h643:rom=16'h6010;
  11'h644:rom=16'h728;
  11'h645:rom=16'h42FF;
  11'h646:rom=16'h2701;
  11'h647:rom=16'hE100;
  11'h648:rom=16'h2FF6;
  11'h649:rom=16'hC020;
  11'h64A:rom=16'h2108;
  11'h64B:rom=16'h6020;
  11'h64C:rom=16'h72A;
  11'h64D:rom=16'h27FF;
  11'h64E:rom=16'h4200;
  11'h64F:rom=16'h3215;
  11'h650:rom=16'h172A;
  11'h651:rom=16'h2FCE;
  11'h652:rom=16'h72A;
  11'h653:rom=16'h42FF;
  11'h654:rom=16'h2701;
  11'h655:rom=16'hE100;
  11'h656:rom=16'h3215;
  11'h657:rom=16'h172A;
  11'h658:rom=16'h2FC3;
  11'h659:rom=16'h170B;
  11'h65A:rom=16'h2FC1;
  11'h65B:rom=16'h170C;
  11'h65C:rom=16'h2FBF;
  11'h65D:rom=16'h3107;
  11'h65E:rom=16'h704;
  11'h65F:rom=16'hC008;
  11'h660:rom=16'h2104;
  11'h661:rom=16'h6008;
  11'h662:rom=16'h171D;
  11'h663:rom=16'h2FC5;
  11'h664:rom=16'h171E;
  11'h665:rom=16'h2FB6;
  11'h666:rom=16'h3107;
  11'h667:rom=16'h705;
  11'h668:rom=16'hC004;
  11'h669:rom=16'h2108;
  11'h66A:rom=16'h6004;
  11'h66B:rom=16'h729;
  11'h66C:rom=16'h27FF;
  11'h66D:rom=16'h4200;
  11'h66E:rom=16'h3215;
  11'h66F:rom=16'h1729;
  11'h670:rom=16'h2FC1;
  11'h671:rom=16'hC008;
  11'h672:rom=16'h2107;
  11'h673:rom=16'h6008;
  11'h674:rom=16'h729;
  11'h675:rom=16'h42FF;
  11'h676:rom=16'h2701;
  11'h677:rom=16'hE100;
  11'h678:rom=16'h2FF6;
  11'h679:rom=16'h3017;
  11'h67A:rom=16'h170F;
  11'h67B:rom=16'hC063;
  11'h67C:rom=16'h2106;
  11'h67D:rom=16'h27EE;
  11'h67E:rom=16'h70E0;
  11'h67F:rom=16'h1E07;
  11'h680:rom=16'h3F80;
  11'h681:rom=16'h2F00;
  11'h682:rom=16'h270D;
  11'h683:rom=16'h710C;
  11'h684:rom=16'hC018;
  11'h685:rom=16'h2F95;
  11'h686:rom=16'h3107;
  11'h687:rom=16'h70F;
  11'h688:rom=16'hC008;
  11'h689:rom=16'h2105;
  11'h68A:rom=16'h6008;
  11'h68B:rom=16'h2701;
  11'h68C:rom=16'h7100;
  11'h68D:rom=16'h2FED;
  11'h68E:rom=16'h2701;
  11'h68F:rom=16'h7101;
  11'h690:rom=16'h2F8B;
  11'h691:rom=16'h2701;
  11'h692:rom=16'h7102;
  11'h693:rom=16'h2F88;
  11'h694:rom=16'h1F11;
  11'h695:rom=16'h1F21;
  11'h696:rom=16'h270D;
  11'h697:rom=16'h2FF9;
  11'h698:rom=16'h2711;
  11'h699:rom=16'h721A;
  11'h69A:rom=16'h228;
  11'h69B:rom=16'h202;
  11'h69C:rom=16'h1E08;
  11'h69D:rom=16'h204;
  11'h69E:rom=16'h1E09;
  11'h69F:rom=16'h1F11;
  11'h6A0:rom=16'h202;
  11'h6A1:rom=16'h216;
  11'h6A2:rom=16'h3018;
  11'h6A3:rom=16'h8000;
  11'h6A4:rom=16'h1202;
  11'h6A5:rom=16'hF11;
  11'h6A6:rom=16'h2708;
  11'h6A7:rom=16'h7000;
  11'h6A8:rom=16'h1E09;
  11'h6A9:rom=16'h270D;
  11'h6AA:rom=16'h2FC9;
  11'h6AB:rom=16'hE00;
  11'h6AC:rom=16'h1E00;
  11'h6AD:rom=16'h2711;
  11'h6AE:rom=16'h721A;
  11'h6AF:rom=16'h229;
  11'h6B0:rom=16'h202;
  11'h6B1:rom=16'h1E08;
  11'h6B2:rom=16'h204;
  11'h6B3:rom=16'h2780;
  11'h6B4:rom=16'h6000;
  11'h6B5:rom=16'h1E09;
  11'h6B6:rom=16'h204;
  11'h6B7:rom=16'h1E09;
  11'h6B8:rom=16'h1F11;
  11'h6B9:rom=16'h202;
  11'h6BA:rom=16'h216;
  11'h6BB:rom=16'h3018;
  11'h6BC:rom=16'h8000;
  11'h6BD:rom=16'h1202;
  11'h6BE:rom=16'hF11;
  11'h6BF:rom=16'h270D;
  11'h6C0:rom=16'h2FC9;
  11'h6C1:rom=16'h204;
  11'h6C2:rom=16'h2780;
  11'h6C3:rom=16'h6000;
  11'h6C4:rom=16'h1E09;
  11'h6C5:rom=16'h2708;
  11'h6C6:rom=16'h7000;
  11'h6C7:rom=16'h1E09;
  11'h6C8:rom=16'h2711;
  11'h6C9:rom=16'h721A;
  11'h6CA:rom=16'h201;
  11'h6CB:rom=16'h9001;
  11'h6CC:rom=16'h1E07;
  11'h6CD:rom=16'h2807;
  11'h6CE:rom=16'h20E;
  11'h6CF:rom=16'h40BF;
  11'h6D0:rom=16'h120E;
  11'h6D1:rom=16'h7000;
  11'h6D2:rom=16'h1E0A;
  11'h6D3:rom=16'h2F0C;
  11'h6D4:rom=16'h1201;
  11'h6D5:rom=16'h20F;
  11'h6D6:rom=16'hC060;
  11'h6D7:rom=16'h2108;
  11'h6D8:rom=16'hE00;
  11'h6D9:rom=16'h2704;
  11'h6DA:rom=16'hC000;
  11'h6DB:rom=16'h29BD;
  11'h6DC:rom=16'h20F;
  11'h6DD:rom=16'hC020;
  11'h6DE:rom=16'h2903;
  11'h6DF:rom=16'h7000;
  11'h6E0:rom=16'h1E09;
  11'h6E1:rom=16'hF21;
  11'h6E2:rom=16'hF11;
  11'h6E3:rom=16'hF00;
  11'h6E4:rom=16'h1F01;
  11'h6E5:rom=16'hF01;
  11'h6E6:rom=16'h1F01;
  11'h6E7:rom=16'hF01;
  11'h6E8:rom=16'h1F01;
  11'h6E9:rom=16'hF01;
  11'h6EA:rom=16'h3F00;
  11'h6EB:rom=16'hF00;
  11'h6EC:rom=16'h21C;
  11'h6ED:rom=16'h7000;
  11'h6EE:rom=16'hC120;
  11'h6EF:rom=16'h2905;
  11'h6F0:rom=16'h7001;
  11'h6F1:rom=16'hC110;
  11'h6F2:rom=16'h2902;
  11'h6F3:rom=16'h9002;
  11'h6F4:rom=16'h1206;
  11'h6F5:rom=16'h2718;
  11'h6F6:rom=16'h7000;
  11'h6F7:rom=16'hC108;
  11'h6F8:rom=16'h2103;
  11'h6F9:rom=16'h2730;
  11'h6FA:rom=16'h6000;
  11'h6FB:rom=16'hF00;
  11'h6FC:rom=16'h270E;
  11'h6FD:rom=16'h2F0F;
  11'h6FE:rom=16'h2F04;
  11'h6FF:rom=16'h2708;
  11'h700:rom=16'h7000;
  11'h701:rom=16'h1E09;
  11'h702:rom=16'hE00;
  11'h703:rom=16'h2701;
  11'h704:rom=16'hC000;
  11'h705:rom=16'h29FA;
  11'h706:rom=16'hF00;
  11'h707:rom=16'hE00;
  11'h708:rom=16'h2702;
  11'h709:rom=16'hC000;
  11'h70A:rom=16'h29FD;
  11'h70B:rom=16'h7000;
  11'h70C:rom=16'h1E09;
  11'h70D:rom=16'hF00;
  11'h70E:rom=16'hF00;
  11'h70F:rom=16'h2711;
  11'h710:rom=16'h702E;
  11'h711:rom=16'h270C;
  11'h712:rom=16'h710A;
  11'h713:rom=16'h1010;
  11'h714:rom=16'h2780;
  11'h715:rom=16'h7100;
  11'h716:rom=16'h1B13;
  11'h717:rom=16'hF00;
  11'h718:rom=16'h00;
  11'h719:rom=16'h3D00;
  11'h71A:rom=16'h393B;
  11'h71B:rom=16'hFF3A;
  11'h71C:rom=16'h00;
  11'h71D:rom=16'h00;
  11'h71E:rom=16'h343C;
  11'h71F:rom=16'h35;
  11'h720:rom=16'h8400;
  11'h721:rom=16'h8281;
  11'h722:rom=16'h1180;
  11'h723:rom=16'h1B;
  11'h724:rom=16'h00;
  11'h725:rom=16'h131A;
  11'h726:rom=16'h1701;
  11'h727:rom=16'h1C;
  11'h728:rom=16'h300;
  11'h729:rom=16'h418;
  11'h72A:rom=16'h1E05;
  11'h72B:rom=16'h1D;
  11'h72C:rom=16'h3300;
  11'h72D:rom=16'h616;
  11'h72E:rom=16'h1214;
  11'h72F:rom=16'h1F;
  11'h730:rom=16'hE00;
  11'h731:rom=16'h802;
  11'h732:rom=16'h1907;
  11'h733:rom=16'h20;
  11'h734:rom=16'h00;
  11'h735:rom=16'hA0D;
  11'h736:rom=16'h2115;
  11'h737:rom=16'h22;
  11'h738:rom=16'h2D00;
  11'h739:rom=16'h90B;
  11'h73A:rom=16'h240F;
  11'h73B:rom=16'h23;
  11'h73C:rom=16'h2E00;
  11'h73D:rom=16'hC2F;
  11'h73E:rom=16'h102B;
  11'h73F:rom=16'h25;
  11'h740:rom=16'h3000;
  11'h741:rom=16'h2C;
  11'h742:rom=16'h2628;
  11'h743:rom=16'h00;
  11'h744:rom=16'h8983;
  11'h745:rom=16'h2931;
  11'h746:rom=16'h2700;
  11'h747:rom=16'h00;
  11'h748:rom=16'h00;
  11'h749:rom=16'h00;
  11'h74A:rom=16'h37;
  11'h74B:rom=16'h32;
  11'h74C:rom=16'h4F00;
  11'h74D:rom=16'h522A;
  11'h74E:rom=16'h55;
  11'h74F:rom=16'h00;
  11'h750:rom=16'h4D4E;
  11'h751:rom=16'h5350;
  11'h752:rom=16'h5654;
  11'h753:rom=16'h4736;
  11'h754:rom=16'h4B00;
  11'h755:rom=16'h4A51;
  11'h756:rom=16'h5749;
  11'h757:rom=16'h38;
  11'h758:rom=16'h00;
  11'h759:rom=16'h00;
  11'h75A:rom=16'h00;
  11'h75B:rom=16'h00;
  11'h75C:rom=16'h00;
  11'h75D:rom=16'h00;
  11'h75E:rom=16'h00;
  11'h75F:rom=16'h00;
  11'h760:rom=16'h8C00;
  11'h761:rom=16'h00;
  11'h762:rom=16'h88;
  11'h763:rom=16'h00;
  11'h764:rom=16'h00;
  11'h765:rom=16'h00;
  11'h766:rom=16'h00;
  11'h767:rom=16'h00;
  11'h768:rom=16'h00;
  11'h769:rom=16'h00;
  11'h76A:rom=16'h00;
  11'h76B:rom=16'h00;
  11'h76C:rom=16'h00;
  11'h76D:rom=16'h00;
  11'h76E:rom=16'h00;
  11'h76F:rom=16'h00;
  11'h770:rom=16'h00;
  11'h771:rom=16'h00;
  11'h772:rom=16'h00;
  11'h773:rom=16'h00;
  11'h774:rom=16'h00;
  11'h775:rom=16'h00;
  11'h776:rom=16'h00;
  11'h777:rom=16'h00;
  11'h778:rom=16'h00;
  11'h779:rom=16'h00;
  11'h77A:rom=16'h00;
  11'h77B:rom=16'h00;
  11'h77C:rom=16'h00;
  11'h77D:rom=16'h48;
  11'h77E:rom=16'h00;
  11'h77F:rom=16'h00;
  11'h780:rom=16'h00;
  11'h781:rom=16'h00;
  11'h782:rom=16'h00;
  11'h783:rom=16'h00;
  11'h784:rom=16'h00;
  11'h785:rom=16'h4C;
  11'h786:rom=16'h00;
  11'h787:rom=16'h00;
  11'h788:rom=16'h00;
  11'h789:rom=16'h00;
  11'h78A:rom=16'h00;
  11'h78B:rom=16'h00;
  11'h78C:rom=16'h00;
  11'h78D:rom=16'h4400;
  11'h78E:rom=16'h42;
  11'h78F:rom=16'h00;
  11'h790:rom=16'h3F3E;
  11'h791:rom=16'h45;
  11'h792:rom=16'h4346;
  11'h793:rom=16'h00;
  11'h794:rom=16'h00;
  11'h795:rom=16'h41;
  11'h796:rom=16'h4000;
  11'h797:rom=16'h00;
  11'h798:rom=16'h3231;
  11'h799:rom=16'h3433;
  11'h79A:rom=16'h3635;
  11'h79B:rom=16'h3837;
  11'h79C:rom=16'h3039;
  11'h79D:rom=16'h5E2D;
  11'h79E:rom=16'h405D;
  11'h79F:rom=16'h5C5B;
  11'h7A0:rom=16'h3A3B;
  11'h7A1:rom=16'h2E2C;
  11'h7A2:rom=16'h5F2F;
  11'h7A3:rom=16'h80D;
  11'h7A4:rom=16'h920;
  11'h7A5:rom=16'h1B1B;
  11'h7A6:rom=16'h13FE;
  11'h7A7:rom=16'h7271;
  11'h7A8:rom=16'h7473;
  11'h7A9:rom=16'h875;
  11'h7AA:rom=16'hE08;
  11'h7AB:rom=16'hB0F;
  11'h7AC:rom=16'h1D1E;
  11'h7AD:rom=16'h1C1F;
  11'h7AE:rom=16'h2F0B;
  11'h7AF:rom=16'h2D2A;
  11'h7B0:rom=16'hD2B;
  11'h7B1:rom=16'h302E;
  11'h7B2:rom=16'h3231;
  11'h7B3:rom=16'h3433;
  11'h7B4:rom=16'h3635;
  11'h7B5:rom=16'h3837;
  11'h7B6:rom=16'hFF39;
  11'h7B7:rom=16'h2221;
  11'h7B8:rom=16'h2423;
  11'h7B9:rom=16'h2625;
  11'h7BA:rom=16'h2827;
  11'h7BB:rom=16'h7E29;
  11'h7BC:rom=16'h603D;
  11'h7BD:rom=16'h607D;
  11'h7BE:rom=16'h7C7B;
  11'h7BF:rom=16'h2A2B;
  11'h7C0:rom=16'h3E3C;
  11'h7C1:rom=16'h5F3F;
  11'h7C2:rom=16'h120D;
  11'h7C3:rom=16'h920;
  11'h7C4:rom=16'h1B1B;
  11'h7C5:rom=16'h3FE;
  11'h7C6:rom=16'h7776;
  11'h7C7:rom=16'h7978;
  11'h7C8:rom=16'h127A;
  11'h7C9:rom=16'hE12;
  11'h7CA:rom=16'hC0F;
  11'h7CB:rom=16'h1D1E;
  11'h7CC:rom=16'h1C1F;
  11'h7CD:rom=16'h2F0C;
  11'h7CE:rom=16'h2D2A;
  11'h7CF:rom=16'hD2B;
  11'h7D0:rom=16'h302E;
  11'h7D1:rom=16'h3231;
  11'h7D2:rom=16'h3433;
  11'h7D3:rom=16'h3635;
  11'h7D4:rom=16'h3837;
  11'h7D5:rom=16'hFF39;
  11'h7D6:rom=16'h3231;
  11'h7D7:rom=16'h3433;
  11'h7D8:rom=16'h3635;
  11'h7D9:rom=16'h3837;
  11'h7DA:rom=16'h3039;
  11'h7DB:rom=16'h1E00;
  11'h7DC:rom=16'h401D;
  11'h7DD:rom=16'h00;
  11'h7DE:rom=16'h00;
  11'h7DF:rom=16'h00;
  11'h7E0:rom=16'h00;
  11'h7E1:rom=16'h0D;
  11'h7E2:rom=16'h00;
  11'h7E3:rom=16'h00;
  11'h7E4:rom=16'h13FE;
  11'h7E5:rom=16'h00;
  11'h7E6:rom=16'h00;
  11'h7E7:rom=16'h00;
  11'h7E8:rom=16'hE00;
  11'h7E9:rom=16'hB0F;
  11'h7EA:rom=16'h1D1E;
  11'h7EB:rom=16'h1C1F;
  11'h7EC:rom=16'h2F0B;
  11'h7ED:rom=16'h2D2A;
  11'h7EE:rom=16'hD2B;
  11'h7EF:rom=16'h302E;
  11'h7F0:rom=16'h3231;
  11'h7F1:rom=16'h3433;
  11'h7F2:rom=16'h3635;
  11'h7F3:rom=16'h3837;
  11'h7F4:rom=16'h39;
  11'h7F5:rom=16'h00;
  11'h7F6:rom=16'h00;
  11'h7F7:rom=16'h00;
  11'h7F8:rom=16'h00;
  11'h7F9:rom=16'h00;
  11'h7FA:rom=16'h00;
  11'h7FB:rom=16'h00;
  11'h7FC:rom=16'h00;
  11'h7FD:rom=16'h00;
  11'h7FE:rom=16'h00;
  11'h7FF:rom=16'h00;
endcase
end
endfunction
/////
always @(posedge CLK)
begin
  DO <= rom(A);
end

endmodule

