// megafunction wizard: %ALTDDIO_BIDIR%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altddio_bidir 

// ============================================================
// File Name: alt_altddio_bidir.v
// Megafunction Name(s):
// 			altddio_bidir
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 350 03/24/2010 SP 2 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2010 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module alt_altddio_bidir (
	aclr,
	datain_h,
	datain_l,
	inclock,
	oe,
	outclock,
	combout,
	dataout_h,
	dataout_l,
	padio);

	input	  aclr;
	input	[0:0]  datain_h;
	input	[0:0]  datain_l;
	input	  inclock;
	input	  oe;
	input	  outclock;
	output	[0:0]  combout;
	output	[0:0]  dataout_h;
	output	[0:0]  dataout_l;
	inout	[0:0]  padio;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri0	  aclr;
	tri1	  oe;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [0:0] sub_wire0;
	wire [0:0] sub_wire1;
	wire [0:0] sub_wire2;
	wire [0:0] dataout_h = sub_wire0[0:0];
	wire [0:0] combout = sub_wire1[0:0];
	wire [0:0] dataout_l = sub_wire2[0:0];

	altddio_bidir	altddio_bidir_component (
				.padio (padio),
				.outclock (outclock),
				.inclock (inclock),
				.oe (oe),
				.datain_h (datain_h),
				.aclr (aclr),
				.datain_l (datain_l),
				.dataout_h (sub_wire0),
				.combout (sub_wire1),
				.dataout_l (sub_wire2),
				.aset (1'b0),
				.dqsundelayedout (),
				.inclocken (1'b1),
				.oe_out (),
				.outclocken (1'b1),
				.sclr (1'b0),
				.sset (1'b0));
	defparam
		altddio_bidir_component.extend_oe_disable = "UNUSED",
		altddio_bidir_component.implement_input_in_lcell = "ON",
		altddio_bidir_component.intended_device_family = "Cyclone II",
		altddio_bidir_component.invert_output = "OFF",
		altddio_bidir_component.lpm_type = "altddio_bidir",
		altddio_bidir_component.oe_reg = "UNUSED",
		altddio_bidir_component.width = 1;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ARESET_MODE NUMERIC "0"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: EXTEND_OE_DISABLE NUMERIC "0"
// Retrieval info: PRIVATE: IMPLEMENT_INPUT_IN_LCELL NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: OE NUMERIC "1"
// Retrieval info: PRIVATE: OE_REG NUMERIC "0"
// Retrieval info: PRIVATE: POWER_UP_HIGH NUMERIC "0"
// Retrieval info: PRIVATE: SRESET_MODE NUMERIC "2"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: USE_COMBOUT NUMERIC "1"
// Retrieval info: PRIVATE: USE_DATAOUT NUMERIC "1"
// Retrieval info: PRIVATE: USE_DQS_UNDELAYOUT NUMERIC "0"
// Retrieval info: PRIVATE: WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: EXTEND_OE_DISABLE STRING "UNUSED"
// Retrieval info: CONSTANT: IMPLEMENT_INPUT_IN_LCELL STRING "ON"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: INVERT_OUTPUT STRING "OFF"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altddio_bidir"
// Retrieval info: CONSTANT: OE_REG STRING "UNUSED"
// Retrieval info: CONSTANT: WIDTH NUMERIC "1"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT GND aclr
// Retrieval info: USED_PORT: combout 0 0 1 0 OUTPUT NODEFVAL combout[0..0]
// Retrieval info: USED_PORT: datain_h 0 0 1 0 INPUT NODEFVAL datain_h[0..0]
// Retrieval info: USED_PORT: datain_l 0 0 1 0 INPUT NODEFVAL datain_l[0..0]
// Retrieval info: USED_PORT: dataout_h 0 0 1 0 OUTPUT NODEFVAL dataout_h[0..0]
// Retrieval info: USED_PORT: dataout_l 0 0 1 0 OUTPUT NODEFVAL dataout_l[0..0]
// Retrieval info: USED_PORT: inclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL inclock
// Retrieval info: USED_PORT: oe 0 0 0 0 INPUT VCC oe
// Retrieval info: USED_PORT: outclock 0 0 0 0 INPUT_CLK_EXT NODEFVAL outclock
// Retrieval info: USED_PORT: padio 0 0 1 0 BIDIR NODEFVAL padio[0..0]
// Retrieval info: CONNECT: @datain_h 0 0 1 0 datain_h 0 0 1 0
// Retrieval info: CONNECT: @datain_l 0 0 1 0 datain_l 0 0 1 0
// Retrieval info: CONNECT: padio 0 0 1 0 @padio 0 0 1 0
// Retrieval info: CONNECT: @outclock 0 0 0 0 outclock 0 0 0 0
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @oe 0 0 0 0 oe 0 0 0 0
// Retrieval info: CONNECT: dataout_h 0 0 1 0 @dataout_h 0 0 1 0
// Retrieval info: CONNECT: dataout_l 0 0 1 0 @dataout_l 0 0 1 0
// Retrieval info: CONNECT: @inclock 0 0 0 0 inclock 0 0 0 0
// Retrieval info: CONNECT: combout 0 0 1 0 @combout 0 0 1 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_altddio_bidir.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_altddio_bidir.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_altddio_bidir.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_altddio_bidir.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_altddio_bidir.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_altddio_bidir_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL alt_altddio_bidir_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
